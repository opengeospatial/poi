"ID"|"Group Number"|"Group Description"
1|"01"|"ACCOMMODATION, EATING AND DRINKING"
2|"02"|"COMMERCIAL SERVICES"
3|"03"|"ATTRACTIONS"
4|"04"|"SPORT AND ENTERTAINMENT"
5|"05"|"EDUCATION AND HEALTH"
6|"06"|"PUBLIC INFRASTRUCTURE"
7|"07"|"MANUFACTURING AND PRODUCTION"
8|"09"|"RETAIL"
9|"10"|"TRANSPORT"
