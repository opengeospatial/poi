PointX Classification Code|Description|First SIC 2003|Second SIC 2003|Third SIC 2003|Fourth SIC 2003|Fifth SIC 2003|Sixth SIC 2003|Seventh SIC 2003|First SIC 2007|Second SIC 2007|Third SIC 2007|Fourth SIC 2007|Fifth SIC 2007|Sixth SIC 2007|Seventh SIC 2007
01010002|Camping, Caravanning, Mobile Homes, Holiday Parks and Centres|5522|5523||||||5530|5520|5590?||||
01010003|Bed and Breakfast and Backpacker Accommodation|5523|||||||5520||||||
01010005|Hostels and Refuges for the Homeless|5523|||||||5590||||||
01010006|Hotels, Motels, Country Houses and Inns|5510|||||||5510||||||
01010007|Self Catering|5523|||||||5520||||||
01010008|Timeshare|5523|||||||5590||||||
01010009|Youth Accommodation|5521|5523||||||5520|5590|||||
01020012|Banqueting and Function Rooms|7020|||||||6820||||||
01020013|Cafes, Snack Bars and Tea Rooms|5530|||||||5610||||||
01020018|Fast Food and Takeaway Outlets|5530|||||||5610||||||
01020019|Fast Food Delivery Services|5530|||||||5610||||||
01020020|Fish and Chip Shops|5530|||||||5610||||||
01020025|Internet Cafes|6420|5530||||||6190|5610|||||
01020034|Pubs, Bars and Inns|5540|||||||5630||||||
01020043|Restaurants|5530|||||||5610||||||
02030044|Metalworkers Including Blacksmiths|2870|2852||||||2599|0162|3311||||
02030045|Building Contractors|4521|4545||||||4120|4339|4399||||
02030046|Construction Completion Services|4545|4534|4532|4542|4525|||4329|4332|4339|3320|4399||
02030047|Construction Plant|2952?|||||||2892?||||||
02030048|Cutting, Drilling and Welding Services|4525|4512|2670|2942|2670|||2562|4313|4221|3311|3312||
02030049|Demolition Services|4511|4550||||||4311|4312|4399||||
02030050|Diving Services|7487?|||||||4291?||||||
02030051|Electrical Contractors|4531|||||||4321|8020?|||||
02030052|Gardening, Landscaping and Tree Surgery Services|0141|7420?||||||8130|0161|||||
02030053|Glaziers|4544|2612|4542?|5246?||||4334|4332|2312?||||
02030054|Painting and Decorating Services|4544|4543||||||4334|4333|||||
02030055|Plasterers|4541|||||||4331||||||
02030056|Plumbing and Heating Services|4533|||||||4322|3311?|||||
02030057|Pool and Court Construction|4523|4545||||||4399||||||
02030058|Restoration and Preservation Services|4545|7470||||||4339|8129|||||
02030059|Road Construction Services|4523|||||||4211||||||
02030060|Roofing and Chimney Services|4522|4525|4531|7470?||||4391|4399|4329|8122?|||
02030778|Fencing and Drystone Walling Services|4525|||||||4399||||||
02030779|Building and Component Suppliers|4543|4542|4525|4534||||4333|4332|4399|4329|||
02040063|Architectural and Building-Related Consultants|7420|4521?||||||7111|7490|||||
02040064|Business-Related Consultants|7414|||||||7022|7490|||||
02040065|Computer Consultants|7222|7210|7230|||||6201|6202|6209|6311|||
02040066|Construction Service Consultants|7420|4532|4533|||||7112|4329|4322||||
02040067|Feng Shui Consultants, Furnishers and Shop Fitters|7487|9305?||||||7410|9609?|||||
02040068|Food Consultants|7430?|8514?|5552?|||||7120?|5629?|8690?||||
02040069|Image Consultants|7414|||||||7021||||||
02040070|Interpretation and Translation Consultants|7485|||||||7430||||||
02040071|Security Consultants|7460|4531||||||7490|8010|8020||||
02040072|Telecommunications Consultants|7487|7420?||||||7490||||||
02040074|Traffic Management and Transport Related Consultants|7487?|6340?|6330?|7420?||||7490?|5229?|7911?||||
02050075|Careers Offices and Armed Forces Recruitment|7450|7522?||||||7810|7820|8422?||||
02050076|Domestic Staff and Home Help|9500|7450||||||9700|7810|7820|8532|8891||
02050077|Driver Agencies|7450|||||||7810|7820|||||
02050078|Employment Agencies|7450|||||||7810|7820|||||
02050079|Modelling and Theatrical Agencies|7487|9272||||||7810|7490|||||
02050081|Nursing Agencies|7450|||||||7810|7820|||||
02060083|Aviation Engineers|7420?|7487?||||||7490?||||||
02060084|Chemical Engineers|7420?|7487?||||||7490?||||||
02060085|Civil Engineers|4521|4523|7420|||||4299|4212|3320|4120|4213|4221|7112
02060086|Electrical and Electronic Engineers|4531|||||||4321||||||
02060087|Hydraulic Engineers|7420|||||||3312|3320?|||||
02060088|Industrial Engineers|7420|||||||3312|3320|||||
02060089|Instrumentation Engineers|7420|||||||3320||||||
02060090|Marine Engineers and Services|6322|7420||||||3315|5222|5020?||||
02060091|Mechanical Engineers|2852|7420||||||3312|2562?|||||
02060092|Pneumatic Engineers|7240|||||||3312|3320|||||
02060093|Precision Engineers|2852|||||||3312|3320|||||
02060094|Structural Engineers|4521|7420||||||4213|4212?|3320?||||
02070095|Agricultural Contractors|0141|7131|4550?|||||7731|7712?|||||
02070096|Aircraft Charters|6220|7123|6210?|||||5110|5121|7735||||
02070098|Catering Services|5552|5551||||||5621|5629|||||
02070100|Contract Cleaning Services|7470|||||||8122|8110|8121|8129|||
02070101|Display and Window Dressers|7440|||||||7311||||||
02070102|Drain and Sewage Clearance|9001|4533?||||||3700|4322?|||||
02070105|Linen Hire and Washroom Services|7470?|9301?||||||8122?|9601?|||||
02070107|Office Services|7133|||||||7733|8219|||||
02070108|Packers|7482|||||||8292||||||
02070109|Pest and Vermin Control|7470|0141?||||||8129|0161?|||||
02080114|Advertising Services|7440|||||||7311|7312|||||
02080115|Artists, Illustrators and Calligraphers|9231|||||||9003||||||
02080116|Computer Security|7222?|7221?||||||6202?|6209?|||||
02080117|Computer Systems Services|7222|7221||||||5821|5829|6201|6209|||
02080118|Concert/Exhibition Organisers and Services|7487|||||||8230||||||
02080119|Database Services|7240|7230||||||6311|6203?|||||
02080120|Desktop Publishing Services|2224|7221?||||||1813|5829|||||
02080121|Electronic and Internet Publishers|7240|||||||5811|5812|5814|5819|5920?||
02080122|Film and Video Services|2232|9211|9220|9213||||1820|5911|5912|5913|||
02080123|General Computer Services|7230|||||||6203|6311|||||
02080124|Internet Services|6420|||||||6190|6312|||||
02080125|Literary Services|7485|9231||||||8211|8219|9003||||
02080126|Mailing and Other Information Services|7240|7485||||||5812|8219|||||
02080127|Marketing Services|7413|||||||7320||||||
02080128|Plate Makers, Print Finishers and Type Setters|2224|||||||1813||||||
02080129|Press and Journalism Services|9240|2224||||||6391|1813|6399|7420|9003||
02080130|Printing and Photocopying Services|7485|2222||||||8219||||||
02080131|Recording Studios and Record Companies|2231|2214||||||1820|5920|||||
02080133|Telephone, Telex and Fax Services|6420|||||||6190||||||
02080134|Television and Radio Services|9220|6420||||||5911|5912|5913|5920|6010|6020|
02090135|Accountants and Auditors|7412|||||||6920||||||
02090137|Auctioneers, Auction Rooms and Valuers|5263|7487||||||4791|8299|||||
02090138|Banks and Building Societies|6512|6511|6523|||||6419|6411|||||
02090140|Currency Conversion and Money Transfers|6713|||||||6612||||||
02090141|Cash Machines|6523?|||||||6499?|9511?|||||
02090142|Cheque Cashing|6713|||||||6619||||||
02090143|Company Registration and Trademarks|7415|7487?||||||6910|7740|||||
02090144|Copyright and Patent|7411|||||||6910|5920|||||
02090145|Credit Reference Agencies|7487|||||||6399|8291|||||
02090146|Debt Collecting Agencies|7487|||||||8291||||||
02090147|Financial Advice Services|6602|6713|6720|||||6530|6520|6619||||
02090148|Fundraising Services|8532|9132|9133|||||8899|9492|9499||||
02090149|Insurers and Support Activities|6601|6603|6720||6523|||6511|6512|6520|6621|6499|6622|6629
02090150|Mortgage and Financial Lenders|6521|6522||||||6491|6492|6499||||
02090151|Pawnbrokers|6522|||||||6492||||||
02090154|Solicitors, Advocates and Notaries Public|7411|||||||6910||||||
02090773|Stocks, Shares and Unit Trusts|6523|6712||||||6430|6499|6612||||
02090795|Commodity Dealers|6523|6711||||||6611|6612|||||
02090796|Franchise and Holding Company Services|6523|7415|7487|||||6420|7010|||||
02090811|PayPoint Locations|7487?|6713?||||||6619||||||
02090829|Pension and Fund Management|6712|6602|6720|||||6630|6430|6530||||
02100103|Hotel Booking Agencies|6330|||||||7990||||||
02100112|Event Ticket Agents and Box Office|9232|6330?||||||7990|7911|||||
02100155|Astrologers, Clairvoyants and Palmists|9305|||||||9609||||||
02100156|Hair and Beauty Services|9302|9304||||||9602|9604|||||
02100158|Cleaning Services|9301|||||||9601||||||
02100160|Customer Service Centres|7486|||||||8220||||||
02100161|CV Writers|9231|9305?||||||9003||||||
02100162|Detective and Investigation Agencies|7460|||||||8030|8010|||||
02100165|Funeral and Associated Services|9303|||||||9603||||||
02100166|Historical Research|9305|9252|9251|||||9609|9102|9101||||
02100167|Headquarters, Administration and Central Offices|7415|||||||7010||||||
02100169|Introduction and Dating Agencies|9305|||||||9609||||||
02100170|Lock, Key and Security Services|2863|5274?||||||2572|8020|4759||||
02100171|Message and Greeting Services|7487?|9234?||||||9001?|8219?|||||
02100173|Motoring Organisations|9133|||||||9499||||||
02100174|Party Organisers|9305?|7487?||||||9609?||||||
02100175|Personalisation|2222?|||||||1812?||||||
02100177|Photographic Services|7481|||||||7420||||||
02100179|Sports Services|9262|||||||9319||||||
02100180|Tattooing and Piercing Services|9305?|||||||9609||||||
02100182|Trophies and Engraving Services|9231|3622|3663|||||9003|3212|3299|9525|||
02100183|Vehicle Cleaning Services|5020|7470?||||||4520|8129?|||||
02100185|Weather Services|7420|||||||7490||||||
02100186|Wedding Services|7481|5552||||||7420|5621|||||
02100188|Window Cleaners|7470|||||||8122||||||
02100774|Musicians, Orchestras and Composers|9231|||||||9001||||||
02100775|Sculptors, Wood Workers and Stone Masons|9231|2670|2051|1411?||||9003|2370|1629|0811|||
02100776|Tailoring and Clothing Alteration|1822|5274||||||1413|9529|||||
02100777|Vehicle Breakdown and Recovery Services|5020|||||||5221||||||
02100818|Sewage Services|9001|||||||3700||||||
02100821|Spas|9304|8514||||||9604|8690|||||
02100822|Slimming Clubs and Services|9133?|1588?||||||9604?|8690?|1086?||||
02100823|Adult Services|9305?|||||||9609?||||||
02100826|Printing on Garments|5274|2222?|1730?|||||1812|1330|||||
02110189|Commercial Property Letting|7020|7031||||||6820|6831|||||
02110190|Property Sales|7031|7011|7012?|||||6831|4110|6810?||||
02110191|Estate and Property Management|7032|7020|7011|||||6820|6832|8110?||||
02110192|Property Letting|7020|||||||6820||||||
02110194|Property Development Services|7011|7012?||||||4110|6810?|||||
02110195|Property Information Services|7420|||||||7111|7112|||||
02120196|Recycling, Reclamation and Disposal|9002|9003||||||3811|3812|3832|8129|||
02120198|Rag Merchants|5157|||||||4677||||||
02120199|Clearance and Salvage Dealers|5157|||||||4677||||||
02120200|Scrap Metal Merchants|3710|5157||||||3832|3831|||||
02120202|Waste Paper Merchants|5157|2111?||||||3811|1711?|4677?||||
02130204|Building Repairs|4525?|4521?|4544?|4545?||||4399?|4334?|4339?||||
02130205|Electrical Equipment Repair and Servicing|7250|5272||||||9511|9521|3312|3313|9512|9522|
02130206|Household Repairs and Restoration|5274|9231|3614?|||||9524|9529|9003?||||
02130207|Industrial Repairs and Servicing|7250|2922||||||3312|3313|4329|3311?|||
02130209|Service Industry Equipment Repairs|5274?|||||||9529?|3312?|3319?||||
02130210|Sports and Leisure Equipment Repair|5274|||||||9529||||||
02130211|Tool Repairs|5274?|2852?||||||3312||||||
02130212|Vehicle Repair, Testing and Servicing|5020|5040|7430|||||4520|3317|4540|7120|||
02130793|Shoe Repairs|5271|||||||9523||||||
02140214|Design Services|7487|7420||||||7410|7111|||||
02140216|Research Services|7310|7320||||||7211|7219|7220||||
02140217|Testing and Analysis Services|7430|||||||7120||||||
02150218|Airlines and Airline Services|6210|6220|6323|||||5110|3316|5121|5223|||
02150219|Animal Transportation|6321|||||||5221||||||
02150221|Container and Storage|6312|7132||||||5210|7739|||||
02150222|Courier, Delivery and Messenger|6412|||||||5320||||||
02150223|Distribution and Haulage|6024|6010|6321|6311|6340|||4941|4920|5221|5224|5229|7490|
02150224|Ferry and Cruise Companies|6110|||||||5010|5020|||||
02150225|Import and Export Services|6340|||||||5229||||||
02150227|Railway Related Services|6010|6321|6021?|||||4910|4920|5221|4931?|||
02150228|Removals and Shipping Agents|6024?|6311?|6340|||||4942|5224?|5229||||
02150230|Taxi Services|6022|||||||4932||||||
02600097|Boat Hiring Services|6110|6120|7122|||||5030|5010|7721|7734|||
02600099|Construction and Tool Hire|7132|7140|4550|||||7732|7739|4399||||
02600104|Leisure Equipment Hirings|7140|||||||7721|7735|||||
02600110|Renting and Leasing of Personal and Household Goods|7140|||||||7729||||||
02600111|Sound, Light and Vision Service and Equipment Hire|7140|||||||7729||||||
02600113|Vehicle Hire and Rental|7110|6023|6022|7121||||7711|4939|7712|7739?|||
02600159|Clothing Hire|7140|9301||||||7729|9601|||||
02600270|Bouncy Castles and Inflatables Hire|9272|||||||9329||||||
03160231|Aquaria and Sea Life Centres|9253|||||||9104||||||
03160232|Bird Reserves, Collections and Sanctuaries|9253|||||||9104||||||
03160233|Butterfly Farms|9253|||||||9104||||||
03160235|Farm Based Attractions|9253?|||||||9104?||||||
03160236|Horticultural Attractions|9253|0141?||||||9104|8130?|||||
03160237|Salmon Ladders|0502|||||||0322||||||
03160239|Zoos and Animal Collections|9253|||||||9104||||||
03170240|Archaeological Sites|9252|||||||9103||||||
03170241|Battlefields|9252|||||||9103||||||
03170244|Historic Buildings Including Castles, Forts and Abbeys|9252|||||||9103||||||
03170245|Historic and Ceremonial Structures|9252|||||||9103||||||
03170246|Historical Ships|9252|||||||9103||||||
03170248|Museums|9252|||||||9102||||||
03170813|Art Galleries|9232|||||||9004||||||
03180252|Commons|9272|9253?||||||9329|9104?|||||
03180253|Country and National Parks|9272?|9253?||||||9329?|9104?|||||
03180254|Picnic Areas|9233?|||||||9321||||||
03180255|Playgrounds|9272|||||||9329||||||
03180814|Municipal Parks and Gardens|0141|||||||8130||||||
03190257|Designated Scenic Features|0000|||||||0000||||||
03190259|Trigonometric Points|7420|||||||7112||||||
03200263|Laseria, Observatories and Planetaria|7310|9232?||||||7219?|9004?|||||
03200264|Model Villages|9234|||||||9321||||||
03200265|Railways (Heritage, Steam and Miniature)|9233|6021|9252|9234||||9329|9103|||||
03200266|Theme and Adventure Parks|9233|||||||9321||||||
03200267|Siteseeing, Tours, Viewing and Visitor Centres|9252|||6110|6120|||9103|9102|||5010|5030|
03200268|Information Centres|6330|||||||7990||||||
03200269|Unspecified and Other Attractions|9252|9272||||||9103|9329|||||
03580803|Ponds|0141?|||||||8130?||||||
03580804|Lakes and Waters|0000|||||||0000||||||
03580805|Lochs and Lochans|0000|||||||0000||||||
03580806|Tarns, Pools and Meres|0000|||||||0000||||||
03580807|Reservoirs|0000|||||||0000||||||
03580808|Settling, Balancing and Silt Ponds|0000|||||||0000||||||
04210271|Children's Activity Centres|9133?|||||||9499?||||||
04210273|Entertainment Services|9234|9231||||||9001|9002|||||
04210274|Firework Related Services|9234|2461||||||9329|2051|||||
04210275|Funfair Services|9233|||||||9321||||||
04210276|Mobile Discos|9234|9231?||||||9329|9001?|||||
04210820|Motorsport Services|9262|||||||9319|9312|||||
04220277|Amusement Parks and Arcades|9271|9272|9233|||||9200|9321|||||
04220278|Bingo Halls|9271|||||||9200||||||
04220279|Bookmakers|9271|||||||9200||||||
04220280|Casinos|9271|||||||9200||||||
04220281|Pools Promoters|9271|||||||9200||||||
04230282|Angling and Sports Fishing|9262|||||||9319||||||
04230283|Combat, Laser and Paintball Games|9272?|||||||9329?||||||
04230284|Hot Air Ballooning|6220?|||||||5110?||||||
04230285|Parachuting and Bungee Jumping|9272?|9262?||||||9329?|9319?|||||
04230286|Paragliding and Hang Gliding|9262?|9272?||||||9319?|9329?|||||
04230287|Watersports|9262|7140?||||||9319|9329|7721?||||
04230321|Riding Schools, Livery Stables and Equestrian Centres|9262|||||||8551|9319?|||||
04230770|Outdoor Pursuit Organisers and Equipment|9262?|9272?|7140?|||||9319?|9329?|7721?||||
04240289|Athletics Facilities|9261|||||||9311||||||
04240290|Bowling Facilities|9261|||||||9311||||||
04240291|Climbing Facilities|9261|||||||9311||||||
04240292|Golf Ranges, Courses, Clubs and Professionals|9261|9262||||||9311|9312|8551?||||
04240293|Gymnasiums, Sports Halls and Leisure Centres|9261|9304||||||9311|9313|||||
04240294|Ice Rinks|9261|||||||9311||||||
04240297|Motorsport Venues|9261|||||||9311||||||
04240298|Racecourses and Greyhound Tracks|9261|||||||9311||||||
04240299|Shooting Facilities|9261|0150||||||9311||||||
04240300|Ski Infrastructure and Aerial Cableways|6021|9261?||||||4939|9311?|||||
04240301|Snooker and Pool Halls|9261|||||||9311||||||
04240302|Sports Grounds, Stadia and Pitches|9261|||||||9311||||||
04240303|Squash Courts|9261|||||||9311||||||
04240304|Swimming Pools|9261|||||||9311||||||
04240305|Tennis Facilities|9261|||||||9311||||||
04240306|Velodromes|9261|||||||9311||||||
04250308|Cinemas|9213|||||||5914||||||
04250311|Discos|5540?|9272?||||||5630?|9329?|||||
04250312|Nightclubs|5540?|9272?||||||5630?|9329?|||||
04250314|Social Clubs|5540|9133||||||5630|9499|||||
04250315|Theatres and Concert Halls|9232|||||||9004|7990?|||||
04250762|Conference and Exhibition Centres|7020|5510?||||||6820|5510?|||||
04250825|Adult Venues|5540?|||||||5630?||||||
05260316|Animal Clipping and Grooming|9305|8520?|0142?|||||9609|7500?|0162?||||
05260317|Dog Training|9305|||||||9609||||||
05260318|Horse Training|9262|9305?||||||9319|9609?|||||
05260319|Kennels and Catteries|9305|||||||9609||||||
05260320|Pet Cemeteries and Crematoria|9303|||||||9603||||||
05260322|Veterinarians and Animal Hospitals|8520|||||||7500||||||
05260323|Veterinary Pharmacies|8520|||||||7500||||||
05270324|Education Authorities|7512|8042?||||||8412|8559?|||||
05270325|Education Services|7512|8042||||||8412|8560|||||
05270326|Examination Boards|7512|||||||8412||||||
05270799|Playing for Success Centres|8042|||||||8560||||||
05270800|Secure Units|8042|||||||8559||||||
05280330|Alternative, Natural and Complementary|8514|9305|9304|||||8690|8551|9604||||
05280333|Foot Related Services|8514|||||||8690||||||
05280335|Dental Technicians|8513|8514||||||8623||||||
05280337|Dieticians and Nutritionists|8514|||||||8690||||||
05280340|Homeopaths|8514|||||||8690||||||
05280342|Midwifery|8514|||||||8690||||||
05280344|Optometrists and Opticians|5248|||||||4778||||||
05280345|Physical Therapy|8514|||||||8690||||||
05280352|Speech Therapists|8514|||||||8690||||||
05280354|Surgeons and Cosmetic Surgeries|8512|||||||8622||||||
05280364|Chemists and Pharmacies|5231|||||||4773||||||
05280365|Clinics and Health Centres|8512|||||||8621||||||
05280367|Dental and Medical Laboratories|8514|3310?|8513?|||||8610|3250?|8623||||
05280368|Dental Surgeries|8513|||||||8623||||||
05280369|Doctors Surgeries|8512|||||||8621||||||
05280370|Hospices|8511|8531?||||||8710||||||
05280371|Hospitals|8511|||||||8610||||||
05280372|Mental Health Centres and Practitioners|8514|||||||8690||||||
05280373|Nursing and Residential Care Homes|8511|8531||||||8710|8720|8790||||
05280780|Accident and Emergency Hospitals|8511|||||||8610||||||
05280809|Parenting and Childcare Services|8532|||||||8899||||||
05280812|Walk-In Centre|8512|8514?||||||8621|8622|8690?||||
05280815|Day and Care Centres|8532|||||||8810||||||
05290106|Medical Equipment Rental and Leasing|7134?|||||||7739?||||||
05290356|Ambulance and Medical Transportation Services|8514|||||||8690||||||
05290357|Blood Transfusion Service|8514|||||||8690||||||
05290358|Counselling and Advice Services|8532|7512|7414?|8514?||||9499|8412|8810|8690?|||
05290359|Health Authorities|7512|||||||8412||||||
05290361|Medical Waste Disposal Services|9002|||||||3822|3821?|||||
05290362|Pregnancy Related Services and Help Centres|8514|||||||8690||||||
05290363|X-Ray Services|8514|||||||8690||||||
05310375|First, Primary and Infant Schools|8010|||||||8520||||||
05310376|Further Education Establishments|8030|||||||8541||||||
05310377|Independent and Preparatory Schools|8021|8010||||||8531|8510|8520||||
05310379|Broad Age Range and Secondary State Schools|8021|||||||8531||||||
05310380|Special Schools and Colleges|8010|8021|8042|8532?||||8520|8531|8891?|8559?|||
05310381|Higher Education Establishments|8030|7310?|7320?|||||8542|7219?|7211?||||
05310382|Unspecified and Other Schools|8042|||||||8559||||||
05310801|Pupil Referral Units|8042|||||||8559||||||
05320384|Ballet and Dance Schools|9234|||||||8552||||||
05320385|Beauty and Hairdressing Schools|8022|||||||8532||||||
05320388|Diving Schools|9262|||||||8532|8551|||||
05320389|Drama Schools|8042|||||||8552||||||
05320390|Driving and Motorcycle Schools|8041|||||||8553||||||
05320391|First Aid Training|8042?|8022?||||||8559|8532?|||||
05320392|Flying Schools|6323|8041||||||5223|8532|8553?||||
05320394|Language Schools|8022|||||||8532||||||
05320395|Martial Arts Instruction|8042|9262?||||||8559|8551?|||||
05320396|Music Teachers and Schools|8022?|8042?||||||8552||||||
05320397|Nursery Schools and Pre and After School Care|8010|8532||||||8510|8891|||||
05320399|Sailing Schools|9262|||||||8553||||||
05320400|Sports and Fitness Coaching|9262|8042?||||||8551|8532?|||||
05320403|Training Providers and Centres|8042|||||||8532|8552|||||
06330404|Armed Services|7522|||||||8422||||||
06330407|Coastal Safety|6322|7524||||||5222|8424|||||
06330408|Consular Services|7521?|7524?||||||8421?|8424?|||||
06330409|Courts, Court Services and Tribunals|7523|||||||8423||||||
06330411|Driving Test Centres|8041?|||||||8553?|8532?|8299?||||
06330412|Embassies and Consulates|9900|7521?||||||9900|8421?|||||
06330414|Fire Brigade Stations|7525|||||||8425||||||
06330415|Central Government|7514|7511|7513|7530|7521|||8411|8413|8430|8899|9101|8421|
06330416|Local Government|7512|7511||||||8412|8411|||||
06330417|Revenue and Customs Offices|7511|||||||8411||||||
06330418|Job Centres|7530|7512||||||8430|8899|||||
06330419|Members of Parliament and Members of European Parliament|7511?|||||||8411?||||||
06330422|Police Stations|7524|||||||8424||||||
06330424|Prisons|7523|||||||8423||||||
06330425|Probation Offices and Police Support Services|7523|7524||||||8423|8424|||||
06330426|Registrars Offices|7511?|||||||8411?||||||
06330429|Social Service Activities|8531|8514|8532|7530?||||8790|8720|8810|8730|8810||
06330431|Tribunals|7411|7523?||||||6910|8423?|||||
06330830|Foreign Country Support Activities|7521?|||||||8421?||||||
06340433|Electrical Features|4013|4012||||||3513|3512|||||
06340435|Fire Safety Features|7525|0202||||||8425|0240|||||
06340437|Gas Features|4022|6030|6312|||||3522|4950|5210||||
06340438|Meteorological Features|7420|||||||7490||||||
06340440|Refuse Disposal Facilities|9002|||||||3821||||||
06340441|Waste Storage, Processing and Disposal|9001|9002||||||3700|3821|||||
06340442|Telecommunications Companies|6420|||||||6110|6120|6130|6190|||
06340443|Telecommunications Features|6420|9220||||||6010|6020|6110|6120|6130|6190|
06340444|Utility Companies and Brokers|4013|4022|4030|4100||||3513|3514|3522|3523|3600||
06340453|Allotments|0112|||||||0113||||||
06340454|Cemeteries and Crematoria|9303|||||||9603||||||
06340455|Drinking Fountains and Water Points|4100?|||||||3600?||||||
06340456|Halls and Community Centres|8532?|7487?|7020?|||||8899?|8230?|||||
06340457|Letter Boxes|6411|||||||5310||||||
06340458|Libraries|9251|||||||9101||||||
06340459|Places of Worship|9131|||||||9491||||||
06340460|Public Telephones|6420|||||||6190||||||
06340461|Public Toilets|9001|||||||3700||||||
06340462|Recycling Centres|3720|9002?||||||3832|3821?|||||
06340802|Wifi Hotspots|6420?|||||||6120?||||||
06350445|Animal Welfare Organisations|9133|||||||9499||||||
06350446|Fan Clubs and Associations|9133|||||||9499||||||
06350447|Sports Clubs and Associations|9262|||||||9312||||||
06350448|Institutes and Professional Organisations|9111|9262|7513|9120|9900|||9411|9420|9900||||
06350449|Political Parties and Related Organisations|9132|||||||9492||||||
06350450|Religious Organisations|9131|||||||9491||||||
06350452|Youth Organisations|9133|||||||9499||||||
06350769|Community Networks and Projects|9133|||||||9499||||||
06350816|Charitable Organisations|9133|||||||9499||||||
06350817|Conservation Organisations|9133|||||||9499||||||
07370464|Baby, Nursery and Playground Equipment|3663|3611?||||||3092|2932|||||
07370465|Beds and Bedding|1740|3615|3611|||||1392|3103|3109||||
07370466|Brushes|3662|||||||3291|2219|||||
07370467|Candles|3663|||||||3299||||||
07370468|Canvas Goods|1740|||||||1392||||||
07370470|Carpets, Flooring, Rugs and Soft Furnishings|1751|5147||||||1393|4673|||||
07370471|Medals, Trophies, Ceremonial and Religious Goods|3622|1740|3663|3150||||3212|1392|3299|2740|||
07370472|China and Glassware|2621|5144?||||||2341|4644?|||||
07370473|Clothing, Components and Accessories|1824|1822|1823|5142||||1413|1414|1419|4642|||
07370474|Cookers and Stoves - Non Electrical|2972|||||||2752||||||
07370475|Cosmetics, Toiletries and Perfumes|2452|2451||||||2042|2041|||||
07370476|Curtains and Blinds|1740|||||||1392||||||
07370477|Cutlery and Tableware|2861|||||||2571||||||
07370478|Disability and Mobility Equipment|3310|3543|4531?|||||2660|3092|3250|2822?|4329?||
07370479|Refrigeration and Freezing Appliances|2971|||||||2751||||||
07370480|Footwear|1930|5142||||||1520|1629|2219|2229|4642||
07370481|Furniture|3611|3612|3613|3614||||3109|3101|3102||||
07370482|Garden Goods|2010|2030|2932|3611|2666|2621?||1610|1623|2830|3109|2369|2341?|
07370483|Giftware|3663?|||||||3299?|2219?|||||
07370485|Hobby, Sports and Pastime Products|3650|3640|1920|3663?||||3240|3230|1512|2899?|||
07370486|Disposable Products|2122|1754?||||||1722||||||
07370487|Jewellery, Gems, Clocks and Watches|3350|3622|3661|5147|5273|||2652|3212|3213|4648|9525||
07370488|Lampshades and Lighting|3150|||||||2740||||||
07370489|Leather Products|1920|1910|5124|1810|1824|||1512|1511|4624|1411|1419||
07370490|Lingerie and Hosiery|1823|1771||||||1414|1431|||||
07370491|Luggage, Bags, Umbrellas and Travel Accessories|1920|3663||||||1512|3299|||||
07370493|Musical Instruments|3630|||||||3220||||||
07370494|Photographic and Optical Equipment|3340|2464|3320?|||||2670|3250|2059|4643|||
07370495|Saunas and Sunbeds|2030|3310?||||||1623|3520?|||||
07370497|Tents, Marquees and Camping Equipment|1740|||||||1392||||||
07370498|Tobacco Products|1600|5125|5135|||||1200|4621|4635||||
07370782|Fireplaces and Mantelpieces|2626?|2670?||||||2320?|2370?|||||
07370785|Conservatories|2811?|||||||2511?||||||
07370790|Bathroom Fixtures, Fittings and Sanitary Equipment|2622|2523|2875|||||2342|2223|2599||||
07380500|Coal Mining|1010|1020||||||0510|0520|0990||||
07380501|Oil and Gas Extraction, Refinery and Product Manufacture|1110|1120|2320|4021||||0610|0620|0910|1920|3521|5221?|5222?
07380502|Ore Mining|1310|1200|1320|||||0710|0721|0729|0990|||
07380503|Peat Extraction|1030|||||||0990||||||
07380504|Sand, Gravel and Clay Extraction and Merchants|1421|1422||||||0812||||||
07380506|Stone Quarrying and Preparation|1411|1412|1413|1450|2670|||0811|0990|2370||||
07380507|Unspecified Quarries Or Mines|1450|1440||||||0899|0990|||||
07390508|Animal Breeders (Not Horses)|0125|||||||0149|0144|||||
07390509|Arable Farming|0111|||||||0111||||||
07390510|Bee Keepers|0125|||||||0149||||||
07390511|Dairy Farming|0121|||||||0141||||||
07390512|Fish and Shellfish|0501|0502|0125|||||0311|0312|0321|0322|||
07390513|Forestry|0201|0202||||||0220|0129|0210|0240|||
07390514|Fruit, Flower and Vegetable Growers|0112|0113|5122|5131||||0113|0124|4622|4631|||
07390515|Hoppers and Silos|6312|||||||5210||||||
07390516|Horse Breeders and Dealers|0122|||||||0143||||||
07390517|Livestock Farming|0123|0122||||||0146|0145|||||
07390518|Mixed Or Unspecified Farming|0130|||||||0150||||||
07390520|Poultry Farming, Equipment and Supplies|0124|||||||0147||||||
07390521|Sheep Dips and Washes|0122?|0142?||||||0145?|0162?|||||
07400522|Alcoholic Drinks|1591|1593|1594|1596|1595|||1101|1102|0121|1103|1104|1105|
07400523|Animal Feeds, Pet Foods, Hay and Straw|1571|1572|5121|5138|3720?|||1091|1092|4621|4638|||
07400524|Baking and Confectionery|1581|1582|1561|1584|5136|||1071|1072|1061|1082|4636||
07400525|Dairy Products|1551|1552|5133|||||1051|1052|4633||||
07400526|Fish, Meat and Poultry Products|1511|1512|1513|1520|5132|5138||1011|1012|1013|1020|1085|4632|4638
07400528|Milling, Refining and Food Additives|1541|1542|1542|1583|1440|1587|5121|1041|1042|1081|1084|4621||
07400529|Non Alcoholic Drinks|1532|1598|4100|||||1032|1107|3600||||
07400530|Catering and Non Specific Food Products|1589|1533||||||1089|1039|||||
07410531|Business Parks and Industrial Estates|0000|||||||0000||||||
07410532|Chimneys|0000|||||||0000||||||
07410533|Conveyors|1010?|1421?|1450?|1411?|1412?|1310?|1320?|0510?|0812?|0899?|0811?|0710?|0729?|
07410534|Energy Production|4011|||||||3511||||||
07410535|Lighting Towers|0000|||||||0000||||||
07410536|Lime Kilns|2652|||||||2352||||||
07410537|Oast Houses|1597|1596?||||||1106|1105?|||||
07410538|Pipelines|6030|||||||4950||||||
07410539|Tanks (Generic)|6312|||||||5210||||||
07410540|Travelling Cranes and Gantries|0000|||||||0000||||||
07410542|Unspecified Works Or Factories|0000|||||||0000||||||
07410543|Water Pumping Stations|4100|6030?|0141?|||||3600|4950?|0161?||||
07420544|Abrasive Products and Grinding Equipment|2681|2451?||||||2391|2041?|||||
07420545|Adhesives and Sealants|2462|||||||2052||||||
07420546|Aeroplanes|3530|||||||3030|2899|||||
07420547|Agricultural Machinery and Goods|2931|2932|5111|5188||||2830|4611|4661||||
07420548|Air and Water Filtration|2923|2924|2971?|||||2825|2829|2751?||||
07420549|Arms and Ammunition|2960|||||||2540||||||
07420550|Bearing, Gear and Drive Elements|2914|||||||2815||||||
07420551|Beekeeping Supplies|2932|||||||2830?||||||
07420553|Bricks, Tiles, Clay and Ceramic Products|2640|2630|2626|2621|2623|2624|2625|2332|2331|2320|2341|2343|2349|
07420555|Cable, Wire and Fibre Optics|2734|2873|2874|3130||||2434|2593|2611|2731|2732|2790|
07420557|Colours, Chemicals and Water Softeners and Supplies|2412|2414|5112|5155|2466|||2012|2014|4612|4675|2059||
07420558|Cleaning Equipment and Supplies|2451|5144||||||2041|4644|||||
07420562|Concrete Products|2651|2661|2663|2664|2665|2666||2351|2361|2363|2364|2365|2369|
07420563|Cooling and Refrigeration|2923|||||||2825||||||
07420564|Electrical Components|3210|5186||||||2611|2612|2733|2790|4652||
07420565|Electrical Motors and Generators|3110|2911||||||2711|2811|||||2530
07420566|Electrical Production and Manipulation Equipment|3120|3140||||||2712|2720|2733|2790|||
07420567|Electronic Equipment|3002|3230|3162|5143|3220|||2620|2640|2651|2630|2790|4643|
07420568|Electronic Media|2465|||||||2680|4652|||||
07420569|Engines|2911|3410|3530|3430||||2811|2910|3030||||
07420571|Fertilisers|2415|1430||||||2015|0891|3821?||||
07420572|Food and Beverage Industry Machinery|2953|||||||2893|2830|||||
07420573|General Construction Supplies|2030|2523|2652|2653|2662|2812|2821/2874|1622|1623|2223|2352|2362|2512|2529/2594
07420574|General Purpose Machinery|2924|2952|5182?|||||2829|2892|4663?||||
07420575|Glass|2611|2613|2615|2612||||2311|2313|2319|2312|||2312
07420576|Horticultural Equipment|2932|2420|5155|||||2830|2020|4675||||
07420577|Industrial Coatings and Finishings|2851|1754|2225|||||2561|1396|1814||||
07420579|Tools Including Machine Shops|2862|2852|2943|2941|2943|2942|5115|2562|2573|2824|2829|2841|2849|4615
07420580|Lifting and Handling Equipment|2922|3420|2932?|||||2822|2920|2830?||||
07420581|Lubricants and Lubricating Equipment|2320|5151|2466|2956?||||1920|4671|2899|2059|||
07420582|Marine Equipment Including Boats and Ships|3511|3512|3320|||||3011|3012|3315|3312|2651||
07420583|Measurement and Inspection Equipment|3320|3162||||||2651||||3250||
07420584|Medical Equipment, Supplies and Pharmaceuticals|2411|2441|2442|3310|5146|||2011|2110|2120|2660|3250|3299|4646
07420585|Metals Manufacturers, Fabricators and Stockholders|2710|2722|2741|2731|2745|2751|2811/2840|2410|2420|2441|2431|2443|2451|2445/2550
07420586|Moulds, Dies and Castings|2862|2943|2956|2951|2751|2753|2754|2573|2849|2841|2891|2451|2453|2454
07420588|Office and Shop Equipment|3001|3612|3611|5185?||||2823|3101|4666?||||
07420589|Ovens and Furnaces|2921|2822?||||||2821|2521?|||||
07420590|Packaging|2040|2522|2871|2872||||1624|2222|2591|2592|||
07420591|Paints, Varnishes and Lacquers|2430|||||||2030||||||
07420594|Pesticides|2420|||||||2020||||||
07420598|Printing Related Machinery|2956|2430|2225?|||||2899|2030|||||
07420599|Published Goods|2211|2222|2221|2223|2212|2213|2215|1811|1814|5811|5812|5813|5814|5819
07420600|Pumps and Compressors|2912|||||||2812|2813|||||
07420601|Radar and Telecommunications Equipment|3230|3162||||||2630||||||
07420602|Road Maintenance Equipment|2952|2320|1450|4523?||||2892|1920|2399|0899|4211?||
07420603|Ropes, Nets and Cordage|1752|||||||1394||||||
07420604|Rubber, Silicones and Plastics|2416|2417|2513|2521|2524|3663||2016|2017|2219|2221|2229|2733|3299
07420605|Seals, Tapes, Taps and Valves|2913|2513||||||2814|2219|2812||||
07420606|Signs|2875|3150|2430|7440|3662?|||2599|2790|2030|5819|3291?||
07420607|Special Purpose Machinery and Equipment|3520|2956|2954|2924?||||3020|2899|2896|2894|2599|2829?|
07420608|Textiles, Fabrics, Silk and Machinery|1711|1712|1713|1715|1717|1730|2954/5141|1310|1320|1330|1391|1396|1399|2894/4641
07420609|Stationery, Stamps, Tags and Labels|2123|3663|2125|5147||||1723|3299|1729|4649|||
07420612|General Manufacturing|3663|2875?|2955?|||||2599|2895|||||
07420613|Vehicle Bodybuilders|3420|||||||2920||||||
07420614|Vehicle Components|3430|2511|3161|2512?|3420?|||2932|2931|2910|2211|2813|2740|
07420615|Vehicles|3410|3541|3542|3543|3550?|||2910|3091|3092||||
07420616|Wood Products Including Charcoal, Paper, Card and Board|2010|2020|2051|2112|2121|2124|2125|1610|1621|1629|1712|1721|1724|1729
07420617|Workwear|1821|1824||||||1412|3299|||||
07420765|Educational Equipment and Supplies|3612|2123|3340?|||||3101|1723|2823|2670|||
07420767|Ice|4030|||||||3530||||||
07420781|Fences, Gates and Railings|2812|2873|2030|||||2512|2593|1623||||
07420783|Access Equipment|2811|2751|2875|4525?||||2511|2599|2451|4399?|||
07420784|Car Ports and Steel Buildings|2811|||||||2511||||||
07420787|Waste Collection, Processing and Disposal Equipment|2523|9001||||||2223|3700|||||
07420788|Glass Fibre Services|2614|||||||2314||||||
07420791|Shelving, Storage, Safes and Vaults|2875|3612||||||2599|3101|||||
09460656|Clothing|5242|5116||||||4771|4616|||||
09460657|Footwear|5243|5116||||||4772|4616|||||
09460659|Jewellery and Fashion Accessories|5248|5273||||||4777|4648|9525||||
09460660|Lingerie and Hosiery|5242|||||||4771||||||
09460797|Baby and Nursery Equipment and Children's Clothes|5242|5248||||||4771|4778|||||
09470661|Bakeries|5224|||||||4724||||||
09470662|Butchers|5222|5132?||||||4722|4632?|||||
09470663|Confectioners|5224|||||||4724||||||
09470665|Delicatessens|5222|5227||||||4722|4729|||||
09470666|Fishmongers|5223|5138||||||4723|4638|||||
09470667|Frozen Foods|5227|5117|5139?|||||4721|4631?|4617?||||
09470668|Green and New Age Goods|5248|5212?||||||4778|4719?|||||
09470669|Grocers, Farm Shops and Pick Your Own|5221|5131|5117|||||4721|4631|4617||||
09470670|Herbs and Spices|5227|5137||||||4729|4637?|||||
09470671|Alcoholic Drinks Including Off Licences and Wholesalers|5225|5134||||||4725|4634|||||
09470672|Organic, Health, Gourmet and Kosher Foods|5227|||||||4729||||||
09470699|Convenience Stores and Independent Supermarkets|5211|5212|5226|5227|5117|||4711|4719|4726|4762|4617||
09470703|Livestock Markets|5111|5123||||||4611|4623|||||
09470705|Markets|5262|||||||4781|4782|4789||||
09470768|Cash and Carry|5190|5117?|5119?|||||4690|4617?|4619?||||
09470798|Tea and Coffee Merchants|5225|5137|5117?|||||4725|4637|4617?||||
09470819|Supermarket Chains|5211|||||||4711||||||
09480674|Books and Maps|5247|5250||||||4761|4779|||||
09480675|Carpets, Rugs, Soft Furnishings and Needlecraft|5248|5241|5116|5141|5147|||4753|4751|4616|4641|4647||
09480676|China and Glassware|5244|5144||||||4759|4644|||||
09480677|Cosmetics, Toiletries, Perfumes and Hairdressing Supplies|5233|5145||||||4775|4645|||||
09480678|Craft Supplies|5248|5247||||||4778|4762|||||
09480679|Cycles and Accessories|5248|5274||||||4764|9529|||||
09480680|Diy and Home Improvement|5246|5154|5113|5153||||4752|4674|4613|4673|4647?||
09480682|Furniture|5244|5147|5185?|||||4759|4647|4665?||||
09480683|Garden Centres and Nurseries|5248|5122||||||4776|4622|||||
09480684|Garden Machinery and Furniture|5246|5244|5147|||||4752|9522|4759|4647|||
09480685|General Household Goods|5244|||||||4759||||||
09480686|Hobby, Sports and Pastime Products|5248|||||||4764|4765|4778||||
09480687|Leather Goods, Luggage and Travel Accessories Including Handbags|5243|5147|5116?|||||4772|4649|4616||||
09480688|Lighting|5244|5143||||||4759|4647|||||
09480689|Music and Video|5245|7140|9251|||||4763|7722|9101||||
09480690|Musical Instruments|5245|||||||4759||||||
09480691|Pets, Supplies and Services|5248|5111?|5138?|||||4776|4611?|4638?||||
09480693|Camping and Caravanning|5248|5010||||||4764|4519|||||
09480694|Travel Agencies|6330|||||||7911|7912|||||
09480700|Department Stores|5212|||||||4719||||||
09480701|Discount Stores|5212|||||||4719||||||
09480704|Mail Order and Catalogue Stores|5261|||||||4791||||||
09480708|Shopping Centres and Retail Parks|0000|||||||0000||||||
09480710|Surplus Goods|5212?|5248?||||||4719?|4778?|||||
09480712|Art and Antiques|5250|9232||||||4779|9004|||||
09480714|Charity Shops|5250|8532||||||4779|8899|||||
09480716|Florists|5248|||||||4776||||||
09480717|Gifts and Cards|5248|||||||4778||||||
09480718|Party Goods and Novelties|5248|||||||4778||||||
09480719|Secondhand Goods|5250|||||||4779||||||
09480720|Computer Supplies|5248|5247?||||||4741|4762?|||||
09480721|Domestic Appliances|5245|||||||4754||||||
09480722|Electrical Goods and Components|5245|||||||4743||||||
09480724|Photographic and Optical Equipment|5248|||||||4778||||||
09480725|Stationery and Office Supplies|5247|5248?||||||4762||||||
09480726|Telephones and Telephone Cards|5248|||||||4742||||||
09480763|Post Offices|6411|||||||5310||||||
09480764|Garages, Garden and Portable Buildings|5248?|||||||4778?||||||
09480766|Fuel Distributors and Suppliers|5112|5151||||||4612|4671|||||
09480824|Adult Shops|5248|||||||4778||||||
09480827|Comics Bookshops|5248?|5247?||||||4778?|4761?|||||
09480828|Computer Shops|5248|5184|3002?|||||4741|4651?|9511?||||
09480831|Potteries|5244|5248||||||4759|4778?|||||
09490695|New Vehicles|5010|5040||||||4511|4519|4540||||
09490696|Secondhand Vehicles|5010|||||||4511|4519|||||
09490697|Vehicle Auctions|5010|||||||4511|4519|||||
09490698|Vehicle Parts and Accessories|5030|||||||4532|4531|||||
10530727|Aeronautical Features|6323|||||||5223||||||
10530728|Airports and Landing Strips|6323|||||||5223||||||
10530729|Helipads|6323|||||||5223||||||
10540730|Bridges|6321?|||||||5221?||||||
10540733|Cattle Grids|0121?|||||||0141?|0142?|||||
10540734|Fords and Level Crossings|6321?|||||||5221?||||||
10540735|Motorway Service Stations|6321?|5530?|5050?|||||5221?|5610?|4730?||||
10540736|Parking|6321|||||||5221||||||
10540737|Petrol and Fuel Stations|5050|||||||4730||||||
10540739|Roadside Telephone Boxes|6321?|||||||5221||||||
10540740|Signalling Facilities|6321|||||||5221||||||
10540742|Tunnels|6321|||||||5221||||||
10540743|Viaducts|6321|||||||5221||||||
10540744|Weighbridges|6321|||||||5221||||||
10550746|Finger Posts, Guide Posts and Cairns|0000|||||||0000||||||
10550747|Footbridges|0000|||||||0000||||||
10550749|Stepping Stones|0000|||||||0000||||||
10550750|Subways|0000|||||||0000||||||
10560751|Aqueducts|6322|||||||5222||||||
10560752|Locks|6322|||||||5222||||||
10560753|Moorings and Unloading Facilities|6322|9262||||||5222|9329|||||
10560754|Rivers and Canal Organisations and Infrastructure|6120|6322||||||5030|5222|||||
10560755|Weirs, Sluices and Dams|6322|||||||5222||||||
10560760|Ferries and Ferry Terminals|6110|6322||||||5010|5020|5222||||
10570731|Bus and Coach Stations, Depots and Companies|6021|6023|6321|||||4939|5221|||||
10570738|Railway Stations, Junctions and Halts|6321|6010?||||||5221||||||
10570756|Tram, Metro and Light Railway Stations and Stops|6021|6321||||||5221|4931?|||||
10570758|Taxi Ranks|6022?|6321?||||||4932?|5221?|||||
10570761|Underground Network Stations|6321|6021?||||||5221|4931?|||||
10570794|London Underground Entrances|6321|6021?||||||5221|4931?|||||
10590732|Bus Stops|6021|||||||4939||||||
10590759|Hail and Ride Zones|6021?|||||||4939?||||||
