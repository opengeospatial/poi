"ID"|"Category Number"|"Category Description"|"Group Number Foreign Key"
1|"01"|"ACCOMMODATION"|"01"
2|"02"|"EATING AND DRINKING"|"01"
3|"03"|"CONSTRUCTION SERVICES"|"02"
4|"04"|"CONSULTANCIES"|"02"
5|"05"|"EMPLOYMENT AND CAREER AGENCIES"|"02"
6|"06"|"ENGINEERING SERVICES"|"02"
7|"07"|"CONTRACT SERVICES"|"02"
8|"08"|"IT, ADVERTISING, MARKETING AND MEDIA SERVICES"|"02"
9|"09"|"LEGAL AND FINANCIAL"|"02"
10|"10"|"PERSONAL, CONSUMER AND OTHER SERVICES"|"02"
11|"11"|"PROPERTY AND DEVELOPMENT SERVICES"|"02"
12|"12"|"RECYCLING SERVICES"|"02"
13|"13"|"REPAIR AND SERVICING"|"02"
14|"14"|"RESEARCH AND DESIGN"|"02"
15|"15"|"TRANSPORT, STORAGE AND DELIVERY"|"02"
16|"16"|"BOTANICAL AND ZOOLOGICAL"|"03"
17|"17"|"HISTORICAL AND CULTURAL"|"03"
18|"18"|"RECREATIONAL"|"03"
19|"19"|"LANDSCAPE FEATURES"|"03"
20|"20"|"TOURISM"|"03"
21|"21"|"SPORT AND ENTERTAINMENT SUPPORT SERVICES"|"04"
22|"22"|"GAMBLING"|"04"
23|"23"|"OUTDOOR PURSUITS"|"04"
24|"24"|"SPORTS COMPLEX"|"04"
25|"25"|"VENUES, STAGE AND SCREEN"|"04"
26|"26"|"ANIMAL WELFARE"|"05"
27|"27"|"EDUCATION SUPPORT SERVICES"|"05"
28|"28"|"HEALTH PRACTITIONERS AND ESTABLISHMENTS"|"05"
29|"29"|"HEALTH SUPPORT SERVICES"|"05"
30|"31"|"PRIMARY, SECONDARY AND TERTIARY EDUCATION"|"05"
31|"32"|"RECREATIONAL AND VOCATIONAL EDUCATION"|"05"
32|"33"|"CENTRAL AND LOCAL GOVERNMENT"|"06"
33|"34"|"INFRASTRUCTURE AND FACILITIES"|"06"
34|"35"|"ORGANISATIONS"|"06"
35|"37"|"CONSUMER PRODUCTS"|"07"
36|"38"|"EXTRACTIVE INDUSTRIES"|"07"
37|"39"|"FARMING"|"07"
38|"40"|"FOODSTUFFS"|"07"
39|"41"|"INDUSTRIAL FEATURES"|"07"
40|"42"|"INDUSTRIAL PRODUCTS"|"07"
41|"46"|"CLOTHING AND ACCESSORIES"|"09"
42|"47"|"FOOD, DRINK AND MULTI ITEM RETAIL"|"09"
43|"48"|"HOUSEHOLD, OFFICE, LEISURE AND GARDEN"|"09"
44|"49"|"MOTORING"|"09"
45|"53"|"AIR"|"10"
46|"54"|"ROAD AND RAIL"|"10"
47|"55"|"WALKING"|"10"
48|"56"|"WATER"|"10"
49|"57"|"PUBLIC TRANSPORT, STATIONS AND INFRASTRUCTURE"|"10"
50|"60"|"HIRE SERVICES"|"02"
51|"58"|"BODIES OF WATER"|"03"
52|"59"|"BUS TRANSPORT"|"10"
