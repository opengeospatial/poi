"Administrative Boundary"|"Area Code"|"Description"
"Aberdeen City"|"UTA"|"Unitary Authority"
"Aberdeenshire"|"UTA"|"Unitary Authority"
"Abertawe - Swansea"|"UTA"|"Unitary Authority"
"Adur District"|"DIS"|"District"
"Allerdale District"|"B"|"Borough"
"Amber Valley District"|"B"|"Borough"
"Angus"|"UTA"|"Unitary Authority"
"Argyll and Bute"|"UTA"|"Unitary Authority"
"Arun District"|"DIS"|"District"
"Ashfield District"|"DIS"|"District"
"Ashford District"|"B"|"Borough"
"Aylesbury Vale District"|"DIS"|"District"
"Babergh District"|"DIS"|"District"
"Barking and Dagenham London Boro"|"LBO"|"London Borough"
"Barnet London Boro"|"LBO"|"London Borough"
"Barnsley District"|"B"|"Borough"
"Barrow-in-Furness District"|"B"|"Borough"
"Basildon District"|"B"|"Borough"
"Basingstoke and Deane District"|"B"|"Borough"
"Bassetlaw District"|"DIS"|"District"
"Bath and North East Somerset"|"UTA"|"Unitary Authority"
"Bedford"|"B"|"Borough"
"Bexley London Boro"|"LBO"|"London Borough"
"Birmingham District"|"B"|"Borough"
"Blaby District"|"DIS"|"District"
"Blackburn with Darwen"|"B"|"Borough"
"Blackpool"|"B"|"Borough"
"Blaenau Gwent - Blaenau Gwent"|"UTA"|"Unitary Authority"
"Bolsover District"|"DIS"|"District"
"Bolton District"|"B"|"Borough"
"Boston District"|"B"|"Borough"
"Bournemouth"|"B"|"Borough"
"Bracknell Forest"|"B"|"Borough"
"Bradford District"|"B"|"Borough"
"Braintree District"|"DIS"|"District"
"Breckland District"|"DIS"|"District"
"Brent London Boro"|"LBO"|"London Borough"
"Brentwood District"|"B"|"Borough"
"Bro Morgannwg - the Vale of Glamorgan"|"UTA"|"Unitary Authority"
"Broadland District"|"DIS"|"District"
"Bromley London Boro"|"LBO"|"London Borough"
"Bromsgrove District"|"DIS"|"District"
"Broxbourne District"|"B"|"Borough"
"Broxtowe District"|"B"|"Borough"
"Burnley District"|"B"|"Borough"
"Bury District"|"B"|"Borough"
"Caerdydd - Cardiff"|"UTA"|"Unitary Authority"
"Caerffili - Caerphilly"|"UTA"|"Unitary Authority"
"Calderdale District"|"B"|"Borough"
"Cambridge District"|"B"|"Borough"
"Camden London Boro"|"LBO"|"London Borough"
"Cannock Chase District"|"DIS"|"District"
"Canterbury District"|"B"|"Borough"
"Carlisle District"|"B"|"Borough"
"Casnewydd - Newport"|"UTA"|"Unitary Authority"
"Castell-nedd Port Talbot - Neath Port Talbot"|"UTA"|"Unitary Authority"
"Castle Point District"|"B"|"Borough"
"Central Bedfordshire"|"UTA"|"Unitary Authority"
"Charnwood District"|"B"|"Borough"
"Chelmsford District"|"B"|"Borough"
"Cheltenham District"|"B"|"Borough"
"Cherwell District"|"DIS"|"District"
"Cheshire East"|"B"|"Borough"
"Cheshire West and Chester"|"B"|"Borough"
"Chesterfield District"|"B"|"Borough"
"Chichester District"|"DIS"|"District"
"Chiltern District"|"DIS"|"District"
"Chorley District"|"B"|"Borough"
"Christchurch District"|"B"|"Borough"
"City and County of the City of London"|"LBO"|"London Borough"
"City of Bristol"|"B"|"Borough"
"City of Derby"|"B"|"Borough"
"City of Edinburgh"|"UTA"|"Unitary Authority"
"City of Kingston upon Hull"|"B"|"Borough"
"City of Leicester"|"B"|"Borough"
"City of Nottingham"|"B"|"Borough"
"City of Peterborough"|"B"|"Borough"
"City of Plymouth"|"B"|"Borough"
"City of Portsmouth"|"B"|"Borough"
"City of Southampton"|"B"|"Borough"
"City of Stoke-on-Trent"|"B"|"Borough"
"City of Westminster London Boro"|"LBO"|"London Borough"
"City of Wolverhampton District"|"B"|"Borough"
"Clackmannanshire"|"UTA"|"Unitary Authority"
"Colchester District"|"B"|"Borough"
"Conwy - Conwy"|"UTA"|"Unitary Authority"
"Copeland District"|"B"|"Borough"
"Corby District"|"B"|"Borough"
"Cornwall"|"UTA"|"Unitary Authority"
"Cotswold District"|"DIS"|"District"
"County Durham"|"UTA"|"Unitary Authority"
"County of Herefordshire"|"UTA"|"Unitary Authority"
"Coventry District"|"B"|"Borough"
"Craven District"|"DIS"|"District"
"Crawley District"|"B"|"Borough"
"Croydon London Boro"|"LBO"|"London Borough"
"Dacorum District"|"B"|"Borough"
"Darlington"|"B"|"Borough"
"Dartford District"|"B"|"Borough"
"Daventry District"|"DIS"|"District"
"Derbyshire Dales District"|"DIS"|"District"
"Doncaster District"|"B"|"Borough"
"Dover District"|"DIS"|"District"
"Dudley District"|"B"|"Borough"
"Dumfries and Galloway"|"UTA"|"Unitary Authority"
"Dundee City"|"UTA"|"Unitary Authority"
"Ealing London Boro"|"LBO"|"London Borough"
"East Ayrshire"|"UTA"|"Unitary Authority"
"East Cambridgeshire District"|"DIS"|"District"
"East Devon District"|"DIS"|"District"
"East Dorset District"|"DIS"|"District"
"East Dunbartonshire"|"UTA"|"Unitary Authority"
"East Hampshire District"|"DIS"|"District"
"East Hertfordshire District"|"DIS"|"District"
"East Lindsey District"|"DIS"|"District"
"East Lothian"|"UTA"|"Unitary Authority"
"East Northamptonshire District"|"DIS"|"District"
"East Renfrewshire"|"UTA"|"Unitary Authority"
"East Riding of Yorkshire"|"UTA"|"Unitary Authority"
"East Staffordshire District"|"B"|"Borough"
"Eastbourne District"|"B"|"Borough"
"Eastleigh District"|"B"|"Borough"
"Eden District"|"DIS"|"District"
"Elmbridge District"|"B"|"Borough"
"Enfield London Boro"|"LBO"|"London Borough"
"Epping Forest District"|"DIS"|"District"
"Epsom and Ewell District"|"B"|"Borough"
"Erewash District"|"B"|"Borough"
"Exeter District"|"B"|"Borough"
"Falkirk"|"UTA"|"Unitary Authority"
"Fareham District"|"B"|"Borough"
"Fenland District"|"DIS"|"District"
"Fife"|"UTA"|"Unitary Authority"
"Forest Heath District"|"DIS"|"District"
"Forest of Dean District"|"DIS"|"District"
"Fylde District"|"B"|"Borough"
"Gateshead District"|"B"|"Borough"
"Gedling District"|"B"|"Borough"
"Glasgow City"|"UTA"|"Unitary Authority"
"Gloucester District"|"B"|"Borough"
"Gosport District"|"B"|"Borough"
"Gravesham District"|"B"|"Borough"
"Great Yarmouth District"|"B"|"Borough"
"Greenwich London Boro"|"LBO"|"London Borough"
"Guildford District"|"B"|"Borough"
"Gwynedd - Gwynedd"|"UTA"|"Unitary Authority"
"Hackney London Boro"|"LBO"|"London Borough"
"Halton"|"B"|"Borough"
"Hambleton District"|"DIS"|"District"
"Hammersmith and Fulham London Boro"|"LBO"|"London Borough"
"Harborough District"|"DIS"|"District"
"Haringey London Boro"|"LBO"|"London Borough"
"Harlow District"|"DIS"|"District"
"Harrogate District"|"B"|"Borough"
"Harrow London Boro"|"LBO"|"London Borough"
"Hart District"|"DIS"|"District"
"Hartlepool"|"B"|"Borough"
"Hastings District"|"B"|"Borough"
"Havant District"|"B"|"Borough"
"Havering London Boro"|"LBO"|"London Borough"
"Hertsmere District"|"B"|"Borough"
"High Peak District"|"B"|"Borough"
"Highland"|"UTA"|"Unitary Authority"
"Hillingdon London Boro"|"LBO"|"London Borough"
"Hinckley and Bosworth District"|"B"|"Borough"
"Horsham District"|"DIS"|"District"
"Hounslow London Boro"|"LBO"|"London Borough"
"Huntingdonshire District"|"DIS"|"District"
"Hyndburn District"|"B"|"Borough"
"Inverclyde"|"UTA"|"Unitary Authority"
"Ipswich District"|"B"|"Borough"
"Isle of Wight"|"UTA"|"Unitary Authority"
"Isles of Scilly"|"UTA"|"Unitary Authority"
"Islington London Boro"|"LBO"|"London Borough"
"Kensington and Chelsea London Boro"|"LBO"|"London Borough"
"Kettering District"|"B"|"Borough"
"King's Lynn and West Norfolk District"|"B"|"Borough"
"Kingston upon Thames London Boro"|"LBO"|"London Borough"
"Kirklees District"|"B"|"Borough"
"Knowsley District"|"B"|"Borough"
"Lambeth London Boro"|"LBO"|"London Borough"
"Lancaster District"|"B"|"Borough"
"Leeds District"|"B"|"Borough"
"Lewes District"|"DIS"|"District"
"Lewisham London Boro"|"LBO"|"London Borough"
"Lichfield District"|"DIS"|"District"
"Lincoln District"|"B"|"Borough"
"Liverpool District"|"B"|"Borough"
"Luton"|"B"|"Borough"
"Maidstone District"|"B"|"Borough"
"Maldon District"|"B"|"Borough"
"Malvern Hills District"|"DIS"|"District"
"Manchester District"|"B"|"Borough"
"Mansfield District"|"DIS"|"District"
"Medway"|"B"|"Borough"
"Melton District"|"B"|"Borough"
"Mendip District"|"DIS"|"District"
"Merthyr Tudful - Merthyr Tydfil"|"UTA"|"Unitary Authority"
"Merton London Boro"|"LBO"|"London Borough"
"Mid Devon District"|"DIS"|"District"
"Mid Suffolk District"|"DIS"|"District"
"Mid Sussex District"|"DIS"|"District"
"Middlesbrough"|"B"|"Borough"
"Midlothian"|"UTA"|"Unitary Authority"
"Milton Keynes"|"B"|"Borough"
"Mole Valley District"|"DIS"|"District"
"Moray"|"UTA"|"Unitary Authority"
"Na h-Eileanan an Iar"|"UTA"|"Unitary Authority"
"New Forest District"|"DIS"|"District"
"Newark and Sherwood District"|"DIS"|"District"
"Newcastle upon Tyne District"|"B"|"Borough"
"Newcastle-under-Lyme District"|"B"|"Borough"
"Newham London Boro"|"LBO"|"London Borough"
"North Ayrshire"|"UTA"|"Unitary Authority"
"North Devon District"|"DIS"|"District"
"North Dorset District"|"DIS"|"District"
"North East Derbyshire District"|"DIS"|"District"
"North East Lincolnshire"|"B"|"Borough"
"North Hertfordshire District"|"DIS"|"District"
"North Kesteven District"|"DIS"|"District"
"North Lanarkshire"|"UTA"|"Unitary Authority"
"North Lincolnshire"|"B"|"Borough"
"North Norfolk District"|"DIS"|"District"
"North Somerset"|"UTA"|"Unitary Authority"
"North Tyneside District"|"B"|"Borough"
"North Warwickshire District"|"B"|"Borough"
"North West Leicestershire District"|"DIS"|"District"
"Northampton District"|"B"|"Borough"
"Northumberland"|"UTA"|"Unitary Authority"
"Norwich District"|"B"|"Borough"
"Nuneaton and Bedworth District"|"B"|"Borough"
"Oadby and Wigston District"|"B"|"Borough"
"Oldham District"|"B"|"Borough"
"Orkney Islands"|"UTA"|"Unitary Authority"
"Oxford District"|"B"|"Borough"
"Pendle District"|"B"|"Borough"
"Pen-y-bont ar Ogwr - Bridgend"|"UTA"|"Unitary Authority"
"Perth and Kinross"|"UTA"|"Unitary Authority"
"Poole"|"B"|"Borough"
"Powys - Powys"|"UTA"|"Unitary Authority"
"Preston District"|"B"|"Borough"
"Purbeck District"|"DIS"|"District"
"Reading"|"B"|"Borough"
"Redbridge London Boro"|"LBO"|"London Borough"
"Redcar and Cleveland"|"B"|"Borough"
"Redditch District"|"B"|"Borough"
"Reigate and Banstead District"|"B"|"Borough"
"Renfrewshire"|"UTA"|"Unitary Authority"
"Rhondda Cynon Taf - Rhondda Cynon Taf"|"UTA"|"Unitary Authority"
"Ribble Valley District"|"B"|"Borough"
"Richmond upon Thames London Boro"|"LBO"|"London Borough"
"Richmondshire District"|"DIS"|"District"
"Rochdale District"|"B"|"Borough"
"Rochford District"|"DIS"|"District"
"Rossendale District"|"B"|"Borough"
"Rother District"|"DIS"|"District"
"Rotherham District"|"B"|"Borough"
"Rugby District"|"B"|"Borough"
"Runnymede District"|"B"|"Borough"
"Rushcliffe District"|"B"|"Borough"
"Rushmoor District"|"B"|"Borough"
"Rutland"|"UTA"|"Unitary Authority"
"Ryedale District"|"DIS"|"District"
"Salford District"|"B"|"Borough"
"Sandwell District"|"B"|"Borough"
"Scarborough District"|"B"|"Borough"
"Scottish Borders"|"UTA"|"Unitary Authority"
"Sedgemoor District"|"DIS"|"District"
"Sefton District"|"B"|"Borough"
"Selby District"|"DIS"|"District"
"Sevenoaks District"|"DIS"|"District"
"Sheffield District"|"B"|"Borough"
"Shepway District"|"DIS"|"District"
"Shetland Islands"|"UTA"|"Unitary Authority"
"Shropshire"|"UTA"|"Unitary Authority"
"Sir Benfro - Pembrokeshire"|"UTA"|"Unitary Authority"
"Sir Ceredigion - Ceredigion"|"UTA"|"Unitary Authority"
"Sir Ddinbych - Denbighshire"|"UTA"|"Unitary Authority"
"Sir Fynwy - Monmouthshire"|"UTA"|"Unitary Authority"
"Sir Gaerfyrddin - Carmarthenshire"|"UTA"|"Unitary Authority"
"Sir y Fflint - Flintshire"|"UTA"|"Unitary Authority"
"Sir Ynys Mon - Isle of Anglesey"|"UTA"|"Unitary Authority"
"Slough"|"B"|"Borough"
"Solihull District"|"B"|"Borough"
"South Ayrshire"|"UTA"|"Unitary Authority"
"South Bucks District"|"DIS"|"District"
"South Cambridgeshire District"|"DIS"|"District"
"South Derbyshire District"|"DIS"|"District"
"South Gloucestershire"|"UTA"|"Unitary Authority"
"South Hams District"|"DIS"|"District"
"South Holland District"|"DIS"|"District"
"South Kesteven District"|"DIS"|"District"
"South Lakeland District"|"DIS"|"District"
"South Lanarkshire"|"UTA"|"Unitary Authority"
"South Norfolk District"|"DIS"|"District"
"South Northamptonshire District"|"DIS"|"District"
"South Oxfordshire District"|"DIS"|"District"
"South Ribble District"|"B"|"Borough"
"South Somerset District"|"DIS"|"District"
"South Staffordshire District"|"DIS"|"District"
"South Tyneside District"|"B"|"Borough"
"Southend-on-Sea"|"B"|"Borough"
"Southwark London Boro"|"LBO"|"London Borough"
"Spelthorne District"|"B"|"Borough"
"St. Albans District"|"B"|"Borough"
"St. Edmundsbury District"|"B"|"Borough"
"St. Helens District"|"B"|"Borough"
"Stafford District"|"B"|"Borough"
"Staffordshire Moorlands District"|"DIS"|"District"
"Stevenage District"|"B"|"Borough"
"Stirling"|"UTA"|"Unitary Authority"
"Stockport District"|"B"|"Borough"
"Stockton-on-Tees"|"B"|"Borough"
"Stratford-on-Avon District"|"DIS"|"District"
"Stroud District"|"DIS"|"District"
"Suffolk Coastal District"|"DIS"|"District"
"Sunderland District"|"B"|"Borough"
"Surrey Heath District"|"B"|"Borough"
"Sutton London Boro"|"LBO"|"London Borough"
"Swale District"|"B"|"Borough"
"Swindon"|"B"|"Borough"
"Tameside District"|"B"|"Borough"
"Tamworth District"|"B"|"Borough"
"Tandridge District"|"DIS"|"District"
"Taunton Deane District"|"B"|"Borough"
"Teignbridge District"|"DIS"|"District"
"Telford and Wrekin"|"B"|"Borough"
"Tendring District"|"DIS"|"District"
"Test Valley District"|"DIS"|"District"
"Tewkesbury District"|"B"|"Borough"
"Thanet District"|"DIS"|"District"
"The City of Brighton and Hove"|"B"|"Borough"
"Three Rivers District"|"DIS"|"District"
"Thurrock"|"B"|"Borough"
"Tonbridge and Malling District"|"B"|"Borough"
"Torbay"|"B"|"Borough"
"Tor-faen - Torfaen"|"UTA"|"Unitary Authority"
"Torridge District"|"DIS"|"District"
"Tower Hamlets London Boro"|"LBO"|"London Borough"
"Trafford District"|"B"|"Borough"
"Tunbridge Wells District"|"B"|"Borough"
"Uttlesford District"|"DIS"|"District"
"Vale of White Horse District"|"DIS"|"District"
"Wakefield District"|"B"|"Borough"
"Walsall District"|"B"|"Borough"
"Waltham Forest London Boro"|"LBO"|"London Borough"
"Wandsworth London Boro"|"LBO"|"London Borough"
"Warrington"|"B"|"Borough"
"Warwick District"|"DIS"|"District"
"Watford District"|"B"|"Borough"
"Waveney District"|"DIS"|"District"
"Waverley District"|"B"|"Borough"
"Wealden District"|"DIS"|"District"
"Wellingborough District"|"B"|"Borough"
"Welwyn Hatfield District"|"B"|"Borough"
"West Berkshire"|"UTA"|"Unitary Authority"
"West Devon District"|"B"|"Borough"
"West Dorset District"|"DIS"|"District"
"West Dunbartonshire"|"UTA"|"Unitary Authority"
"West Lancashire District"|"B"|"Borough"
"West Lindsey District"|"DIS"|"District"
"West Lothian"|"UTA"|"Unitary Authority"
"West Oxfordshire District"|"DIS"|"District"
"West Somerset District"|"DIS"|"District"
"Weymouth and Portland District"|"B"|"Borough"
"Wigan District"|"B"|"Borough"
"Wiltshire"|"UTA"|"Unitary Authority"
"Winchester District"|"B"|"Borough"
"Windsor and Maidenhead"|"B"|"Borough"
"Wirral District"|"B"|"Borough"
"Woking District"|"B"|"Borough"
"Wokingham"|"B"|"Borough"
"Worcester District"|"B"|"Borough"
"Worthing District"|"B"|"Borough"
"Wrecsam - Wrexham"|"UTA"|"Unitary Authority"
"Wychavon District"|"DIS"|"District"
"Wycombe District"|"DIS"|"District"
"Wyre District"|"B"|"Borough"
"Wyre Forest District"|"DIS"|"District"
"York"|"B"|"Borough"
