Keyword or phrase|Group|Category1|Category2|Category3|Class1|Class2|Class3|Class4|Class5|comment
Abattoir|||||526|||||
Accommodation agencies|||||192|||||
Accounting, book-keeping and tax services|||||135|147||||
Acupuncture|||||330|||||
Adult education||31|32||376|403||||
Advertising, public relations and marketing agencies|||||114|||||
After school clubs|||||397|452||||
Agricultural colleges|||||403|||||
Agriculture raw materials|||||571|547||||
Air transport||15|53||96|218|728|||
Air transport equipment hire|||||96|392|284|||
Aircrafts / spacecrafts|||||615|546||||probably too generic or for spacecraft not applicable?
Airports|||||728|||||
Alcoholic drinks||47|||522|671||||
Amusement arcades|||||277|||||
Animal boarding premises|||||319|||||
Animal feed mills|||||523|245||||
Animal feeding stuffs||40|39||523|691|520|515||
Animal grooming|||||316|321||||
Animal sanctuaries|||||239|||||
Animal training|||||317|318||||
Antique shops|||||712|719||||
Arable farming|||||509|||||
Architecture / surveying|||||63|195||||
Aromatherapy|||||330|677||||
Art and craft shops|||||712|676||||
Art and illustrations|||||115|712||||
Art studios|||||115|775||||
Auctioneering|||||137|||||
Baby equipment shops|||||797|464||||
Bakery / confectionary|||||661|663|524|572||
Banks|||||138|||||
Beauty salons|||||156|||||
Beauty shops|||||677|||||
Bed and breakfasts - licensed|||||3|||||Not a specific mapping
Bed and breakfasts - non licensed|||||3|||||Not a specific mapping
Bed sits|||||192|||||
Betting shops|||||279|||||
Beverages|||||798|671|522|529|13|Not a specific term and could be mapped to many classes
Bicycle shops|||||679|||||
Bingo halls|||||278|||||
Bird removal|||||416|446||||Not specific assumed environmental health and RSPB type activity?
Boat building (and components)|||||582|686|90|||
Boat hire|||||97|267||||
Boat yard|||||582|753|90|||
Book shops|||||674|827||||
Books|||||674|599||||
Bowling alleys|||||290|||||
Bowls clubs|||||290|||||
Bread and flour||47|||528|524||||
Brewery|||||522|||||
Builders' merchant shops|||||680|779||||
Builders' merchants services||3|48|||||||
Building contracting||3|||45|771|46|||
Building materials|||||680|553|573|504||Not very specific and can be taken to be in a lot of classes
Building societies|||||138|||||
Bureau de changes|||||140|||||
Bus / coach transport|||||731|732|759|267|113|
Business and management consultancies|||||64|||||
Butchery|||||526|662||||
Cafes - licensed|||||13|||||not specific breakdown
Cafes - non-licensed|||||13|||||not specific breakdown
Cakes / pastries / biscuits / pies|||||524|661||||
Camping shops|||||693|||||
Campsites and caravan parks|||||2|||||
Canteens||||||||||Not really held
Car trading - private address|||||696|695||||
Caravan showrooms|||||693|||||
Card / gift shops|||||676|||||
Cargo handling and storage||15|||225|223|221|||
Carpet laying|||||675|46||||not specifically identified
Carpets|||||675|470||||
Cash and carry|||||768|||||
Casinos and gambling clubs|||||280|||||
Cat breeding|||||508|||||
Cattle farming|||||517|511|518|||
Ceramics / non-metal mineral products|||||553|504||||not particularly specific
Charitable organisations|||||816|450||||
Charity shops|||||714|||||
Cheese making|||||525|||||
Chemists / pharmacies|||||364|||||
Childminding and nanny services|||||397|76||||
Children's homes|||||429|||||
Chiropody and podiatry|||||333|||||
Chiropractics and osteopathy|||||345|||||
Cinemas|||||308|||||
Civil engineering||3|||85|||||
Clothes shops|||||656|||||
Clothing and shoes|||||473|480||||Manufacturing and Production version
Clothing and shoes|||||656|657||||Wholesale version
Clothing, textiles and shoe designing|||||214|||||
Coach and bus hire|||||113|||||
Coal|||||500|766||||
Coal merchants' shops|||||766|||||
Coffin making shops|||||165|||||
Coke / petroleum products / nuclear fuel||38|||500|501||||
Computer / office equipment shops|||||828|720|725|||
Computer related activities||4|8||65|117|116|828|720|Very broad could also include class 0100 etc
Confectionary|||||663|||||Wholesale has none retail is shown
Confectionary / chocolates / sugar|||||524|||||Manufacturing
Conference centres|||||762|||||
Construction products||42|||786|||||Manufacturing
Consulting||4|3||64|||||Various classes across groups specified
Consumer credit broking|||||150|||||
Cosmetics|||||677|||||Manufacture
Cosmetics|||||677|||||Wholesale
Counselling services|||||358|||||
Courier services|||||222|||||
Dairy (milk) rounds|||||222|||||unsure if this is included?
Dairy farming|||||511|||||
Dairy produce|||||665|699||||wholesale of food
Dairy products|||||525|||||Manufacturing of food
Data processing and database activities|||||119|||||
Day nurseries|||||397|||||
Debt recovery services|||||146|||||
Delicatessen|||||665|||||
Dental services|||||368|335|584|||
Department stores|||||700|||||
Distribution|||||223|||||
Doctor's surgeries|||||369|||||
Dog breeding|||||508|||||
Do-it-yourself shops|||||680|||||
Domestic chemicals, rubber and plastics|||||558|604||||Manufacturing of
Domestic electrical equipment|||||479|||||Manufacturing of
Double glazing shops|||||680|204||||
Driving schools|||||390|||||
Dry cleaning and launderette services|||||158|||||
Ear / body piercing services|||||180|||||
Editorial and literary services|||||125|||||
Egg packing|||||108|||||unsure if actually in this class or not
Egg producing|||||526|520||||
Egg stalls||47|||520|669||||Retail of
Eggs|||||520|526||||Wholesale
Electrical appliance shops|||||720|||||
Electrical goods|||||720|||||
Electrical installation|||||51|86||||
Electrical machinery / equipment|||||565|479|564|||Manufacturing of
Electricity supply|||||444|433|534|||
Electrology|||||156|330||||
Embalming services|||||165|||||Taxidermists?
Emergency locksmith shops|||||170|||||not specifically emergency
Engineering|||||88|85||||potentially many more
Estate agents' services||9|||190|192||||
Events and exhibitions services|||||118|||||
Extra-territorial organizations||35|||446|816|445|817||Not for profit organisations
Fairgrounds|||||266|||||Amusement parks is 277, Funfair services 275
Farm and agricultural supplies|||||547|95||||
Farm shops|||||669|||||
Farmers market|||||669|672||||not specifically farmers markets
Fertilisers|||||571|||||
Film and video production|||||122|||||
Financial advise / consulting|||||147|150||||
Financial intermediation services|||||448|147||||
Fish / seafoods|||||526|||||wholesale
Fish and fish products|||||512|526||||manufacturing
Fishing and fish farming|||||512|||||
Fishing tackle shops|||||686|||||
Fishmongers|||||666|||||
Fitness and sports centres|||||293|||||
Floor and wall covering|||||54|46||||construction and building services
Florist shops and floral displays|||||716|||||
Flowers|||||683|716|514|||wholesale
Flying / gliding clubs|||||392|286||||
Food haulage (non-live)|||||223|||||
Food importing|||||225|||||
Food packing|||||590|108||||
Forestry (including logging)|||||513|52||||
Forestry consulting|||||513|||||
Frozen food centres|||||667|||||
Fruit and vegetables|||||669|||||wholesale
Fruit farming / orchards|||||514|||||
Fruit packing|||||108|590||||
Fruits and vegetables|||||514|||||manufacturing
Funeral director services|||||165|||||
Funeral services|||||165|||||
Furniture (non-upholstered)|||||682|684||||wholesale
Furniture and upholstery|||||481|588||||Manufacture
Furniture and upholstery|||||682|684||||Retail
Furniture and upholstery shops|||||682|684||||
Game propagation|||||520|508||||Game covers both birds, rabbits, deer etc
Garage - new motor vehicles|||||695|||||
Garage - second-hand motor vehicles|||||696|||||
Garden centres|||||683|||||
General stores|||||699|819||||
Glass / glazing products|||||575|||||manufacturing
Glazing||3|||53|204||||
Goat farming|||||508|517||||possibly even 518?
Golf clubs|||||292|||||
Graphic designing|||||115|214||||
Greengrocer shops|||||669|||||
Grounds maintenance and landscaping|||||52|||||
Guesthouses|||||3|||||
Gunsmith shops|||||686|||||
Haberdashers' shops|||||675|||||
Hackney carriage licensee|||||230|||||
Hackney carriage operators|||||230|||||
Hairdressing salons|||||156|||||
Hairdressing services|||||156|385|677|||
Hardware|||||786|||||
Hardware consultancies|||||65|||||
Hardware shops|||||680|||||
Haulage - non-food|||||223|222||||
Health authorities registered nursing homes|||||373|||||not necessarily registered
Health food shops|||||672|669||||
Herbal shops|||||670|672||||
Higher education institutions||32|||376|||||
Holiday cottages / chalets|||||7|||||
Home catering|||||7|76||||unsure of exact context for this!
Homeopathy|||||340|||||
Horse keeping|||||516|321||||
Horticultural supplies|||||576|683|684|||Class 0576 is down as manufacture but is more
Horticulture / nurseries|||||514|683||||
Hospital kitchens||||||||||not really catered for!
Hospitals|||||371|||||
Hostels|||||5|9||||
Hotels|||||6|3||||
Household / personal goods repair shops|||||206|793|204|211||
Household and leisure equipment||37||||||||Manufacture
Household goods||48|||680|||||Wholesale
Hunt kennels|||||319|||||not believed to be held as such
Industrial cleaning services|||||100|||||
Insurance services|||||149|||||
Interior designing|||||214|||||
Ironmongers shops|||||680|||||
Jewellery|||||487|||||Manufacture
Jewellery shops|||||659|||||Retail
Joinery|||||46|573||||
Knackers' yard|||||526|||||
Landlord tenancy|||||192|||||not specifically held
Lawnmowers and garden machinery|||||684|683|547|||Retail
Legal services|||||154|||||
Leisure centres|||||293|||||
Libraries|||||458|||||
Lighting equipment / furniture shops||48|||688|682|680|||
Liquid fuels / minerals / chemicals||38|||766|536||||Wholesale
Live animals|||||508|520|703|||Wholesale
Livestock auctioneering|||||508|703|137|||Not sure if in 137 and whether others are really relevant
Livestock haulage|||||223|||||
Locksmith shops|||||170|||||
Luncheon clubs||||||||||not catered for?
Machinery||42||||||||Manufacturing
Machinery / equipment rental|||||99|107|111|789||Business service
Machines / equipment||42||||||||Wholesale
Mail order businesses|||||704|||||
Malting|||||537|528||||
Management of holding companies|||||143|||||add in lcc 1855 poss class 150 and 773
Market gardens|||||514|453||||453 is not necessarily a direct mapping
Market stalls|||||705|||||not specifically in
Market stalls (non-food)|||||705|||||not specifically in
Masseurs / masseuse services|||||345|||||Not specifically in this class as it is more medical
Meat and meat products|||||526|662||||Manufacturing - NB no linkage for producers
Meat and meat products|||||526|662||||Wholesale - NB no linkage for producers
Meat packing|||||526|108||||
Mechanical engineering||42|||91|||||Manufacturing
Meditation and Hypnotherapy|||||372|||||
Members' only organisations||35|||314|448||||
Metals|||||585|||||Manufacturing
Milk|||||511|||||Wholesale
Milk bottling|||||511|||||
Milk distributing|||||223|||||
Mixed farming|||||518|||||
Mobile phones and telecommunications|||||442|443|133|72||
Mobile shops||||||||||Not in PointX as no fixed location
Modelling agencies|||||79|||||
Money lending services|||||150|151||||
Motor parts and accessories retail|||||698|||||
Motor vehicle servicing / garage services|||||212|777||||
Motor vehicles / parts / accessories|||||615|547||||Manufacturing
Motorcycles / bicycles|||||615|||||Manufacturing
Motorvehicles and accessories|||||615|547||||Wholesale
Museum / gallery shops|||||712|676||||Retail
Museums / galleries|||||248|813||||
Music / recording studios|||||131|||||
Musical instrument shops|||||690|||||
News agencies (food outlet)|||||699|||||no differentiation between food and non
News agencies (non-food)|||||699|||||no differentiation between food and non
Nightclubs|||||312|825||||825 is more likely to be strip clubs and Pole dancing venues
Non-agricultural raw materials||38|42||524|528|553|557||Wholesale - not very specific!
Non-alcoholic beverages|||||529|||||Wholesale
Non-commercial stables|||||321|||||what is meant by non-commercial? Most here are likely to be
Non-domestic chemicals|||||557|||||Manufacturing
Non-domestic electrical equipment||42||||||||Manufacturing
Non-food importing|||||225|||||
Non-food packing|||||108|590||||
Non-licensed riding stables|||||321|||||
Nursing agencies|||||81|76||||
Nursing homes|||||373|370||||
Off-licences|||||671|||||
Optometric services|||||344|||||
Organic farming||39||||||||not differentiated
Other foods||40|39|||||||Manufacture
Other foods||47|40|39||||||Wholesale
Other land transport||54||||||||other to what???!!
Other livestock farming||39|||517|508||||
Other transport equipment||42||||||||unsure what this means!
Outside catering|||||98|||||
Paint shops|||||680|676||||
Painting and decorating services|||||54|204||||only lcc 2345 from class 204
Pastoral farming|||||517|518||||
Pawn broking shops|||||151|||||
Pensions|||||829|147||||
Performing arts||25|||273|315||||
Personal protective equipment|||||617|||||
Personal training, aerobics, yoga and dance services|||||400|384|330|||
Personnel and recruitment services||5|||78|75||||
Pet food|||||691|523||||Wholesale
Pet shops|||||691|||||
Petrol station (without shop)|||||737|||||records without a corresponding entry in class 699
Petrol station with shops|||||737|||||will have a corresponding entry in class 699
Petroleum and gas supply|||||444|766|501|538||
Pharmaceutical goods|||||584|364||||Wholesale
Photography|||||177|115||||service: 115 much less so
Photography shops|||||724|177||||177 much less so in this context
Physiotherapy|||||345|||||
Piano tuning services|||||210|||||
Picture framing|||||177|206||||service
Picture framing shops|||||177|206||||retail
Pig farming|||||517|518||||518 much less so
Plant hire and tool rental|||||99|||||
Plastering|||||46|45||||45 much less so
Playgroups|||||397|||||
Plumbing and heating services|||||56|||||service could also include 46 and 51 at a stretch
Ports / docks|||||753|97||||97 less so
Post office|||||763|||||
Poultry farming|||||520|||||
Poultry products|||||526|||||
Printing / publishing|||||599|129|121|||129 and even 115 less so
Printing, paper and packaging|||||590|599|616|||Manufacturing Primarily 590.
Private hire licensee|||||113|230||||rental
Private hire operators|||||113|230||||rental
Private investigation and surveillance services|||||162|||||
Private schools|||||379|376||||376 much less so
Property letting / sale / purchase|||||190|192|195|||
Public houses and bars|||||34|||||
Quarantine premises||||||||||Not specifically identified as such
Quarrying / extraction||38|||506|504||||all in category applicable
Radio and television|||||134|443||||
Rail transport||54|||227|265||||
Railway / tramway / rolling stock|||||615|227||||neither of suggestions are really specific
Real estate auctioneering|||||137|||||
Recorded media|||||568|||||Manufacture
Recorded music / video / games shops|||||689|686||||Retail
Recycling||12||||||||
Reflexology|||||345|||||
Regulatory bodies|||||448|415||||
Removal services|||||223|||||
Research organisations / special interest groups|||||216|448|446|173||
Residential clubs|||||8|||||unsure exactly what this is!
Residential homes|||||373|||||
Residential homes and care workers|||||373|370|429|81|76|Drop off in likely relevancy
Restaurants - licensed|||||43|||||
Restaurants - non-licensed|||||43|||||
Riding / livery establishments|||||321|516|318|||
Roadside catering|||||18|13|43|||not really applicable in "mobile" sense
Roofing / thatching contracting|||||60|||||
Saddlery|||||485|||||
School kitchens||||||||||not catered for!
School meals production||||||||||not catered for!
Schools / colleges|||||379|376||||
Second hand-shops|||||719|714||||
Secretarial / admin / personal assistant services|||||78|||||
Security services|||||71|170|791|||not as in MI5 etc!
Self-catering accommodation|||||7|||||
Sewage works|||||441|||||
Sex shops|||||824|||||
Sheep farming|||||517|518|521|||
Shoe repair / key cutting shops|||||793|170||||
Shoe shops|||||657|||||
Shopfittings|||||46|588|67|||
Skip hire|||||99|||||
Social work|||||429|||||
Software consultancies|||||117|65|116|||
Solicitors' services|||||154|||||
Soups / condiments / seasonings|||||530|528||||Manufacturing
Sports grounds|||||302|289|293|||
Sports shops|||||686|770||||
Static alarm consulting|||||71|||||unsure exactly what this is?
Stationery|||||609|725||||Wholesale
Stationery shops|||||725|||||
Stock brokerage|||||773|||||
Sun beds / solariums|||||156|293||||class 293 much less so
Supermarkets|||||819|699||||
Swimming pools and water sports|||||304|287||||
Takeaways|||||18|13|43|||classes 13 and 43 less so
Tattooing|||||180|||||
Taxis and minicabs|||||230|||||
Telephone shops (including mobiles)|||||726|||||
Television / electrical repair service|||||720|||||
Textiles (not clothing)|||||608|675|225|||Wholesale
Textiles and leather (not clothing)||37|42||608|470||||Manufacturing
Theatres|||||315|||||
Ticket booking agencies|||||694|307||||
Timber management|||||513|52||||
Tobacco and tobacco products|||||498|||||Manufacturing
Tobacco products|||||699|||||Wholesale
Tobacco shops|||||699|||||Retail
Toy shops|||||686|||||
Toys / games / sports equipment|||||686|485||||Wholesale NB Distributors so not overlap with retail as normally
Toys / games / sports equipment|||||485|||||Manufacturing
Translation services|||||70|||||
Transport agencies||15|||448|74||||unsure of exact meaning in this context
Travel agencies / tour operator companies|||||694|267||||
Tree maintenance|||||52|513||||
Trichology|||||156|||||
Tyre / exhaust fitting|||||212|||||
Vegetable growing|||||514|453||||
Vehicle alarm consulting|||||71|||||
Vehicle rental|||||113|||||
Vehicles auctioneering|||||697|||||
Veterinary services|||||322|323||||
Video / computer game rental|||||689|||||mainly retail but rental included
Vocational Courses||32|||403|||||
Waste / Scrap||12||||||||
Watch repair shops|||||659|||||possibly also in 487
Water / soft drinks|||||529|444||||Manufacturing
Water services and supplies|||||444|543|455|529||
Water transport||56|15||760|224||||
Web developing|||||117|65|124|||
Wedding and party services|||||186|174||||
Weigh and save shops||47||||||||unsure which specific class will be in as not held as such
Wine / spirits / other beverages|||||671|522|225|||Wholesale
Wood|||||513|616||||Manufacturing
Wood shops|||||766|775|616|||not really retail?
Wool shops|||||675|||||
Zoos|||||239|235||||235 might not exist 231 for Aquaria
