"ID"|"Class Number"|"Classification Description"|"Category Number Foreign Key"
1|"0002"|"CAMPING, CARAVANNING, MOBILE HOMES, HOLIDAY PARKS AND CENTRES"|"01"
2|"0003"|"BED AND BREAKFAST AND BACKPACKER ACCOMMODATION"|"01"
3|"0005"|"HOSTELS AND REFUGES FOR THE HOMELESS"|"01"
4|"0006"|"HOTELS, MOTELS, COUNTRY HOUSES AND INNS"|"01"
5|"0007"|"SELF CATERING"|"01"
6|"0008"|"TIMESHARE"|"01"
7|"0009"|"YOUTH ACCOMMODATION"|"01"
8|"0012"|"BANQUETING AND FUNCTION ROOMS"|"02"
9|"0013"|"CAFES, SNACK BARS AND TEA ROOMS"|"02"
10|"0018"|"FAST FOOD AND TAKEAWAY OUTLETS"|"02"
11|"0019"|"FAST FOOD DELIVERY SERVICES"|"02"
12|"0020"|"FISH AND CHIP SHOPS"|"02"
13|"0025"|"INTERNET CAFES"|"02"
14|"0034"|"PUBS, BARS AND INNS"|"02"
15|"0043"|"RESTAURANTS"|"02"
16|"0044"|"METALWORKERS INCLUDING BLACKSMITHS"|"03"
17|"0045"|"BUILDING CONTRACTORS"|"03"
18|"0046"|"CONSTRUCTION COMPLETION SERVICES"|"03"
19|"0047"|"CONSTRUCTION PLANT"|"03"
20|"0048"|"CUTTING, DRILLING  AND WELDING SERVICES"|"03"
21|"0049"|"DEMOLITION SERVICES"|"03"
22|"0050"|"DIVING SERVICES"|"03"
23|"0051"|"ELECTRICAL CONTRACTORS"|"03"
24|"0052"|"GARDENING, LANDSCAPING AND TREE SURGERY SERVICES"|"03"
25|"0053"|"GLAZIERS"|"03"
26|"0054"|"PAINTING AND DECORATING SERVICES"|"03"
27|"0055"|"PLASTERERS"|"03"
28|"0056"|"PLUMBING AND HEATING SERVICES"|"03"
29|"0057"|"POOL AND COURT CONSTRUCTION"|"03"
30|"0058"|"RESTORATION AND PRESERVATION SERVICES"|"03"
31|"0059"|"ROAD CONSTRUCTION SERVICES"|"03"
32|"0060"|"ROOFING AND CHIMNEY SERVICES"|"03"
33|"0778"|"FENCING AND DRYSTONE WALLING SERVICES"|"03"
34|"0779"|"BUILDING AND COMPONENT SUPPLIERS"|"03"
35|"0063"|"ARCHITECTURAL AND BUILDING RELATED CONSULTANTS"|"04"
36|"0064"|"BUSINESS RELATED CONSULTANTS"|"04"
37|"0065"|"COMPUTER CONSULTANTS"|"04"
38|"0066"|"CONSTRUCTION SERVICE CONSULTANTS"|"04"
39|"0067"|"FENG SHUI CONSULTANTS, FURNISHERS AND SHOP FITTERS"|"04"
40|"0068"|"FOOD CONSULTANTS"|"04"
41|"0069"|"IMAGE CONSULTANTS"|"04"
42|"0070"|"INTERPRETATION AND TRANSLATION CONSULTANTS"|"04"
43|"0071"|"SECURITY CONSULTANTS"|"04"
44|"0072"|"TELECOMMUNICATIONS CONSULTANTS"|"04"
45|"0074"|"TRAFFIC MANAGEMENT AND TRANSPORT RELATED CONSULTANTS"|"04"
46|"0075"|"CAREERS OFFICES AND ARMED FORCES RECRUITMENT"|"05"
47|"0076"|"DOMESTIC STAFF AND HOME HELP"|"05"
48|"0077"|"DRIVER AGENCIES"|"05"
49|"0078"|"EMPLOYMENT AGENCIES"|"05"
50|"0079"|"MODELLING AND THEATRICAL AGENCIES"|"05"
51|"0081"|"NURSING AGENCIES"|"05"
52|"0083"|"AVIATION ENGINEERS"|"06"
53|"0084"|"CHEMICAL ENGINEERS"|"06"
54|"0085"|"CIVIL ENGINEERS"|"06"
55|"0086"|"ELECTRICAL AND ELECTRONIC ENGINEERS"|"06"
56|"0087"|"HYDRAULIC ENGINEERS"|"06"
57|"0088"|"INDUSTRIAL ENGINEERS"|"06"
58|"0089"|"INSTRUMENTATION ENGINEERS"|"06"
59|"0090"|"MARINE ENGINEERS AND SERVICES"|"06"
60|"0091"|"MECHANICAL ENGINEERS"|"06"
61|"0092"|"PNEUMATIC ENGINEERS"|"06"
62|"0093"|"PRECISION ENGINEERS"|"06"
63|"0094"|"STRUCTURAL ENGINEERS"|"06"
64|"0095"|"AGRICULTURAL CONTRACTORS"|"07"
65|"0096"|"AIRCRAFT CHARTERS"|"07"
66|"0098"|"CATERING SERVICES"|"07"
67|"0100"|"CONTRACT CLEANING SERVICES"|"07"
68|"0101"|"DISPLAY AND WINDOW DRESSERS"|"07"
69|"0102"|"DRAIN AND SEWAGE CLEARANCE"|"07"
70|"0105"|"LINEN HIRE AND WASHROOM SERVICES"|"07"
71|"0107"|"OFFICE SERVICES"|"07"
72|"0108"|"PACKERS"|"07"
73|"0109"|"PEST AND VERMIN CONTROL"|"07"
74|"0114"|"ADVERTISING SERVICES"|"08"
75|"0115"|"ARTISTS, ILLUSTRATORS AND CALLIGRAPHERS"|"08"
76|"0116"|"COMPUTER SECURITY"|"08"
77|"0117"|"COMPUTER SYSTEMS SERVICES"|"08"
78|"0118"|"CONCERT/EXHIBITION ORGANISERS AND SERVICES"|"08"
79|"0119"|"DATABASE SERVICES"|"08"
80|"0120"|"DESKTOP PUBLISHING SERVICES"|"08"
81|"0121"|"ELECTRONIC AND INTERNET PUBLISHERS"|"08"
82|"0122"|"FILM AND VIDEO SERVICES"|"08"
83|"0123"|"GENERAL COMPUTER SERVICES"|"08"
84|"0124"|"INTERNET SERVICES"|"08"
85|"0125"|"LITERARY SERVICES"|"08"
86|"0126"|"MAILING AND OTHER INFORMATION SERVICES"|"08"
87|"0127"|"MARKETING SERVICES"|"08"
88|"0128"|"PLATE MAKERS, PRINT FINISHERS AND TYPE SETTERS"|"08"
89|"0129"|"PRESS AND JOURNALISM SERVICES"|"08"
90|"0130"|"PRINTING AND PHOTOCOPYING SERVICES"|"08"
91|"0131"|"RECORDING STUDIOS AND RECORD COMPANIES"|"08"
92|"0133"|"TELEPHONE, TELEX AND FAX SERVICES"|"08"
93|"0134"|"TELEVISION AND RADIO SERVICES"|"08"
94|"0135"|"ACCOUNTANTS AND AUDITORS"|"09"
95|"0137"|"AUCTIONEERS, AUCTION ROOMS AND VALUERS"|"09"
96|"0138"|"BANKS AND BUILDING SOCIETIES"|"09"
97|"0140"|"CURRENCY CONVERSION AND MONEY TRANSFERS"|"09"
98|"0141"|"CASH MACHINES"|"09"
99|"0142"|"CHEQUE CASHING"|"09"
100|"0143"|"COMPANY REGISTRATION AND TRADEMARKS"|"09"
101|"0144"|"COPYRIGHT AND PATENT"|"09"
102|"0145"|"CREDIT REFERENCE AGENCIES"|"09"
103|"0146"|"DEBT COLLECTING AGENCIES"|"09"
104|"0147"|"FINANCIAL ADVICE SERVICES"|"09"
105|"0148"|"FUNDRAISING SERVICES"|"09"
106|"0149"|"INSURERS AND SUPPORT ACTIVITIES"|"09"
107|"0150"|"MORTGAGE AND FINANCIAL LENDERS"|"09"
108|"0151"|"PAWNBROKERS"|"09"
109|"0154"|"SOLICITORS, ADVOCATES AND NOTARIES PUBLIC"|"09"
110|"0773"|"STOCKS, SHARES AND UNIT TRUSTS"|"09"
111|"0795"|"COMMODITY DEALERS"|"09"
112|"0796"|"FRANCHISE AND HOLDING COMPANY SERVICES"|"09"
113|"0811"|"PAYPOINT LOCATIONS"|"09"
114|"0829"|"PENSION AND FUND MANAGEMENT"|"09"
115|"0103"|"HOTEL BOOKING AGENCIES"|"10"
116|"0112"|"EVENT TICKET AGENTS AND BOX OFFICE"|"10"
117|"0155"|"ASTROLOGERS, CLAIRVOYANTS AND PALMISTS"|"10"
118|"0156"|"HAIR AND BEAUTY SERVICES"|"10"
119|"0158"|"CLEANING SERVICES"|"10"
120|"0160"|"CUSTOMER SERVICE CENTRES"|"10"
121|"0161"|"CV WRITERS"|"10"
122|"0162"|"DETECTIVE AND INVESTIGATION AGENCIES"|"10"
123|"0165"|"FUNERAL AND ASSOCIATED SERVICES"|"10"
124|"0166"|"HISTORICAL RESEARCH"|"10"
125|"0167"|"HEADQUARTERS, ADMINISTRATION AND CENTRAL OFFICES"|"10"
126|"0169"|"INTRODUCTION AND DATING AGENCIES"|"10"
127|"0170"|"LOCK, KEY AND SECURITY SERVICES"|"10"
128|"0171"|"MESSAGE AND GREETING SERVICES"|"10"
129|"0173"|"MOTORING ORGANISATIONS"|"10"
130|"0174"|"PARTY ORGANISERS"|"10"
131|"0175"|"PERSONALISATION"|"10"
132|"0177"|"PHOTOGRAPHIC SERVICES"|"10"
133|"0179"|"SPORTS SERVICES"|"10"
134|"0180"|"TATTOOING AND PIERCING SERVICES"|"10"
135|"0182"|"TROPHIES AND ENGRAVING SERVICES"|"10"
136|"0183"|"VEHICLE CLEANING SERVICES"|"10"
137|"0185"|"WEATHER SERVICES"|"10"
138|"0186"|"WEDDING SERVICES"|"10"
139|"0188"|"WINDOW CLEANERS"|"10"
140|"0774"|"MUSICIANS, ORCHESTRAS AND COMPOSERS"|"10"
141|"0775"|"SCULPTORS, WOOD WORKERS AND STONE MASONS"|"10"
142|"0776"|"TAILORING AND CLOTHING ALTERATION"|"10"
143|"0777"|"VEHICLE BREAKDOWN AND RECOVERY SERVICES"|"10"
144|"0818"|"SEWAGE SERVICES"|"10"
145|"0821"|"SPAS"|"10"
146|"0822"|"SLIMMING CLUBS AND SERVICES"|"10"
147|"0823"|"ADULT SERVICES"|"10"
148|"0826"|"PRINTING ON GARMENTS"|"10"
149|"0189"|"COMMERCIAL PROPERTY LETTING"|"11"
150|"0190"|"PROPERTY SALES"|"11"
151|"0191"|"ESTATE AND PROPERTY MANAGEMENT"|"11"
152|"0192"|"PROPERTY LETTING"|"11"
153|"0194"|"PROPERTY DEVELOPMENT SERVICES"|"11"
154|"0195"|"PROPERTY INFORMATION SERVICES"|"11"
155|"0196"|"RECYCLING, RECLAMATION AND DISPOSAL"|"12"
156|"0198"|"RAG MERCHANTS"|"12"
157|"0199"|"CLEARANCE AND SALVAGE DEALERS"|"12"
158|"0200"|"SCRAP METAL DEALERS AND BREAKERS YARDS"|"12"
159|"0202"|"WASTE PAPER MERCHANTS"|"12"
160|"0204"|"BUILDING REPAIRS"|"13"
161|"0205"|"ELECTRICAL EQUIPMENT REPAIR AND SERVICING"|"13"
162|"0206"|"HOUSEHOLD REPAIRS AND RESTORATION"|"13"
163|"0207"|"INDUSTRIAL REPAIRS AND SERVICING"|"13"
164|"0209"|"SERVICE INDUSTRY EQUIPMENT REPAIRS"|"13"
165|"0210"|"SPORTS AND LEISURE EQUIPMENT REPAIR"|"13"
166|"0211"|"TOOL REPAIRS"|"13"
167|"0212"|"VEHICLE REPAIR, TESTING AND SERVICING"|"13"
168|"0793"|"SHOE REPAIRS"|"13"
169|"0214"|"DESIGN SERVICES"|"14"
170|"0216"|"RESEARCH SERVICES"|"14"
171|"0217"|"TESTING AND ANALYSIS SERVICES"|"14"
172|"0218"|"AIRLINES AND AIRLINE SERVICES"|"15"
173|"0219"|"ANIMAL TRANSPORTATION"|"15"
174|"0221"|"CONTAINER AND STORAGE"|"15"
175|"0222"|"COURIER, DELIVERY AND MESSENGER"|"15"
176|"0223"|"DISTRIBUTION AND HAULAGE"|"15"
177|"0224"|"FERRY AND CRUISE COMPANIES"|"15"
178|"0225"|"IMPORT AND EXPORT SERVICES"|"15"
179|"0227"|"RAILWAY RELATED SERVICES"|"15"
180|"0228"|"REMOVALS AND SHIPPING AGENTS"|"15"
181|"0230"|"TAXI SERVICES"|"15"
182|"0097"|"BOAT HIRING SERVICES"|"60"
183|"0099"|"CONSTRUCTION AND TOOL HIRE"|"60"
184|"0104"|"LEISURE EQUIPMENT HIRINGS"|"60"
185|"0110"|"RENTING AND LEASING OF PERSONAL AND HOUSEHOLD GOODS"|"60"
186|"0111"|"SOUND, LIGHT AND VISION SERVICE AND EQUIPMENT HIRE"|"60"
187|"0113"|"VEHICLE HIRE AND RENTAL"|"60"
188|"0159"|"CLOTHING HIRE"|"60"
189|"0270"|"BOUNCY CASTLES AND INFLATABLES HIRE"|"60"
190|"0231"|"AQUARIA AND SEA LIFE CENTRES"|"16"
191|"0232"|"BIRD RESERVES, COLLECTIONS AND SANCTUARIES"|"16"
192|"0233"|"BUTTERFLY FARMS"|"16"
193|"0235"|"FARM BASED ATTRACTIONS"|"16"
194|"0236"|"HORTICULTURAL ATTRACTIONS"|"16"
195|"0237"|"SALMON LADDERS"|"16"
196|"0239"|"ZOOS AND ANIMAL COLLECTIONS"|"16"
197|"0240"|"ARCHAEOLOGICAL SITES"|"17"
198|"0241"|"BATTLEFIELDS"|"17"
199|"0244"|"HISTORIC BUILDINGS INCLUDING CASTLES, FORTS AND ABBEYS"|"17"
200|"0245"|"HISTORIC AND CEREMONIAL STRUCTURES"|"17"
201|"0246"|"HISTORICAL SHIPS"|"17"
202|"0248"|"MUSEUMS"|"17"
203|"0813"|"ART GALLERIES"|"17"
204|"0252"|"COMMONS"|"18"
205|"0253"|"COUNTRY AND NATIONAL PARKS"|"18"
206|"0254"|"PICNIC AREAS"|"18"
207|"0255"|"PLAYGROUNDS"|"18"
208|"0814"|"MUNICIPAL PARKS AND GARDENS"|"18"
209|"0257"|"DESIGNATED SCENIC FEATURES"|"19"
210|"0259"|"TRIGONOMETRIC POINTS"|"19"
211|"0263"|"LASERIA, OBSERVATORIES AND PLANETARIA"|"20"
212|"0264"|"MODEL VILLAGES"|"20"
213|"0265"|"RAILWAYS (HERITAGE, STEAM AND MINIATURE)"|"20"
214|"0266"|"THEME AND ADVENTURE PARKS"|"20"
215|"0267"|"SITESEEING, TOURS, VIEWING AND VISITOR CENTRES"|"20"
216|"0268"|"INFORMATION CENTRES"|"20"
217|"0269"|"UNSPECIFIED AND OTHER ATTRACTIONS"|"20"
218|"0803"|"PONDS"|"58"
219|"0804"|"LAKES AND WATERS"|"58"
220|"0805"|"LOCHS AND LOCHANS"|"58"
221|"0806"|"TARNS, POOLS AND MERES"|"58"
222|"0807"|"RESERVOIRS"|"58"
223|"0808"|"SETTLING, BALANCING AND SILT PONDS"|"58"
224|"0271"|"CHILDREN'S ACTIVITY CENTRES"|"21"
225|"0273"|"ENTERTAINMENT SERVICES"|"21"
226|"0274"|"FIREWORK RELATED SERVICES"|"21"
227|"0275"|"FUNFAIR SERVICES"|"21"
228|"0276"|"MOBILE DISCOS"|"21"
229|"0820"|"MOTORSPORT SERVICES"|"21"
230|"0277"|"AMUSEMENT PARKS AND ARCADES"|"22"
231|"0278"|"BINGO HALLS"|"22"
232|"0279"|"BOOKMAKERS"|"22"
233|"0280"|"CASINOS"|"22"
234|"0281"|"POOLS PROMOTERS"|"22"
235|"0282"|"ANGLING AND SPORTS FISHING"|"23"
236|"0283"|"COMBAT, LASER AND PAINTBALL GAMES"|"23"
237|"0284"|"HOT AIR BALLOONING"|"23"
238|"0285"|"PARACHUTING AND BUNGEE JUMPING"|"23"
239|"0286"|"PARAGLIDING AND HANG GLIDING"|"23"
240|"0287"|"WATERSPORTS"|"23"
241|"0321"|"RIDING SCHOOLS, LIVERY STABLES AND EQUESTRIAN CENTRES"|"23"
242|"0770"|"OUTDOOR PURSUIT ORGANISERS AND EQUIPMENT"|"23"
243|"0289"|"ATHLETICS FACILITIES"|"24"
244|"0290"|"BOWLING FACILITIES"|"24"
245|"0291"|"CLIMBING FACILITIES"|"24"
246|"0292"|"GOLF RANGES, COURSES, CLUBS AND PROFESSIONALS"|"24"
247|"0293"|"GYMNASIUMS, SPORTS HALLS AND LEISURE CENTRES"|"24"
248|"0294"|"ICE RINKS"|"24"
249|"0297"|"MOTORSPORT VENUES"|"24"
250|"0298"|"RACECOURSES AND GREYHOUND TRACKS"|"24"
251|"0299"|"SHOOTING FACILITIES"|"24"
252|"0300"|"SKI INFRASTRUCTURE AND AERIAL CABLEWAYS"|"24"
253|"0301"|"SNOOKER AND POOL HALLS"|"24"
254|"0302"|"SPORTS GROUNDS, STADIA AND PITCHES"|"24"
255|"0303"|"SQUASH COURTS"|"24"
256|"0304"|"SWIMMING POOLS"|"24"
257|"0305"|"TENNIS FACILITIES"|"24"
258|"0306"|"VELODROMES"|"24"
259|"0308"|"CINEMAS"|"25"
260|"0311"|"DISCOS"|"25"
261|"0312"|"NIGHTCLUBS"|"25"
262|"0314"|"SOCIAL CLUBS"|"25"
263|"0315"|"THEATRES AND CONCERT HALLS"|"25"
264|"0762"|"CONFERENCE AND EXHIBITION CENTRES"|"25"
265|"0825"|"ADULT VENUES"|"25"
266|"0316"|"ANIMAL CLIPPING AND GROOMING"|"26"
267|"0317"|"DOG TRAINING"|"26"
268|"0318"|"HORSE TRAINING"|"26"
269|"0319"|"KENNELS AND CATTERIES"|"26"
270|"0320"|"PET CEMETERIES AND CREMATORIA"|"26"
271|"0322"|"VETERINARIANS AND ANIMAL HOSPITALS"|"26"
272|"0323"|"VETERINARY PHARMACIES"|"26"
273|"0324"|"EDUCATION AUTHORITIES"|"27"
274|"0325"|"EDUCATION SERVICES"|"27"
275|"0326"|"EXAMINATION BOARDS"|"27"
276|"0799"|"PLAYING FOR SUCCESS CENTRES"|"27"
277|"0800"|"SECURE UNITS"|"27"
278|"0330"|"ALTERNATIVE, NATURAL AND COMPLEMENTARY"|"28"
279|"0333"|"FOOT RELATED SERVICES"|"28"
280|"0335"|"DENTAL TECHNICIANS"|"28"
281|"0337"|"DIETICIANS AND NUTRITIONISTS"|"28"
282|"0340"|"HOMEOPATHS"|"28"
283|"0342"|"MIDWIFERY"|"28"
284|"0344"|"OPTOMETRISTS AND OPTICIANS"|"28"
285|"0345"|"PHYSICAL THERAPY"|"28"
286|"0352"|"SPEECH THERAPISTS"|"28"
287|"0354"|"SURGEONS AND COSMETIC SURGERIES"|"28"
288|"0364"|"CHEMISTS AND PHARMACIES"|"28"
289|"0365"|"CLINICS AND HEALTH CENTRES"|"28"
290|"0367"|"DENTAL AND MEDICAL LABORATORIES"|"28"
291|"0368"|"DENTAL SURGERIES"|"28"
292|"0369"|"DOCTORS SURGERIES"|"28"
293|"0370"|"HOSPICES"|"28"
294|"0371"|"HOSPITALS"|"28"
295|"0372"|"MENTAL HEALTH CENTRES AND PRACTITIONERS"|"28"
296|"0373"|"NURSING AND RESIDENTIAL CARE HOMES"|"28"
297|"0780"|"ACCIDENT AND EMERGENCY HOSPITALS"|"28"
298|"0809"|"PARENTING AND CHILDCARE SERVICES"|"28"
299|"0812"|"WALK-IN CENTRE"|"28"
300|"0815"|"DAY AND CARE CENTRES"|"28"
301|"0106"|"MEDICAL EQUIPMENT RENTAL AND LEASING"|"29"
302|"0356"|"AMBULANCE AND MEDICAL TRANSPORTATION SERVICES"|"29"
303|"0357"|"BLOOD TRANSFUSION SERVICE"|"29"
304|"0358"|"COUNSELLING AND ADVICE SERVICES"|"29"
305|"0359"|"HEALTH AUTHORITIES"|"29"
306|"0361"|"MEDICAL WASTE DISPOSAL SERVICES"|"29"
307|"0362"|"PREGNANCY RELATED SERVICES AND HELP CENTRES"|"29"
308|"0363"|"X-RAY SERVICES"|"29"
309|"0375"|"FIRST, PRIMARY AND INFANT SCHOOLS"|"31"
310|"0376"|"FURTHER EDUCATION ESTABLISHMENTS"|"31"
311|"0377"|"INDEPENDENT AND PREPARATORY SCHOOLS"|"31"
312|"0379"|"BROAD AGE RANGE AND SECONDARY STATE SCHOOLS"|"31"
313|"0380"|"SPECIAL SCHOOLS AND COLLEGES"|"31"
314|"0381"|"HIGHER EDUCATION ESTABLISHMENTS"|"31"
315|"0382"|"UNSPECIFIED AND OTHER SCHOOLS"|"31"
316|"0801"|"PUPIL REFERRAL UNITS"|"31"
317|"0384"|"BALLET AND DANCE SCHOOLS"|"32"
318|"0385"|"BEAUTY AND HAIRDRESSING SCHOOLS"|"32"
319|"0388"|"DIVING SCHOOLS"|"32"
320|"0389"|"DRAMA SCHOOLS"|"32"
321|"0390"|"DRIVING AND MOTORCYCLE SCHOOLS"|"32"
322|"0391"|"FIRST AID TRAINING"|"32"
323|"0392"|"FLYING SCHOOLS"|"32"
324|"0394"|"LANGUAGE SCHOOLS"|"32"
325|"0395"|"MARTIAL ARTS INSTRUCTION"|"32"
326|"0396"|"MUSIC TEACHERS AND SCHOOLS"|"32"
327|"0397"|"NURSERY SCHOOLS AND PRE AND AFTER SCHOOL CARE"|"32"
328|"0399"|"SAILING SCHOOLS"|"32"
329|"0400"|"SPORTS AND FITNESS COACHING"|"32"
330|"0403"|"TRAINING PROVIDERS AND CENTRES"|"32"
331|"0404"|"ARMED SERVICES"|"33"
332|"0407"|"COASTAL SAFETY"|"33"
333|"0408"|"CONSULAR SERVICES"|"33"
334|"0409"|"COURTS, COURT SERVICES AND TRIBUNALS"|"33"
335|"0411"|"DRIVING TEST CENTRES"|"33"
336|"0412"|"EMBASSIES AND CONSULATES"|"33"
337|"0414"|"FIRE BRIGADE STATIONS"|"33"
338|"0415"|"CENTRAL GOVERNMENT"|"33"
339|"0416"|"LOCAL GOVERNMENT"|"33"
340|"0417"|"REVENUE AND CUSTOMS OFFICES"|"33"
341|"0418"|"JOB CENTRES"|"33"
342|"0419"|"MEMBERS OF PARLIAMENT AND MEMBERS OF EUROPEAN PARLIAMENT"|"33"
343|"0422"|"POLICE STATIONS"|"33"
344|"0424"|"PRISONS"|"33"
345|"0425"|"PROBATION OFFICES AND POLICE SUPPORT SERVICES"|"33"
346|"0426"|"REGISTRARS OFFICES"|"33"
347|"0429"|"SOCIAL SERVICE ACTIVITIES"|"33"
348|"0431"|"TRIBUNALS"|"33"
349|"0830"|"FOREIGN COUNTRY SUPPORT ACTIVITIES"|"33"
350|"0433"|"ELECTRICAL FEATURES"|"34"
351|"0435"|"FIRE SAFETY FEATURES"|"34"
352|"0437"|"GAS FEATURES"|"34"
353|"0438"|"METEOROLOGICAL FEATURES"|"34"
354|"0440"|"REFUSE DISPOSAL FACILITIES"|"34"
355|"0441"|"WASTE STORAGE, PROCESSING AND DISPOSAL"|"34"
356|"0442"|"TELECOMMUNICATIONS COMPANIES"|"34"
357|"0443"|"TELECOMMUNICATIONS FEATURES"|"34"
358|"0444"|"UTILITY COMPANIES AND BROKERS"|"34"
359|"0453"|"ALLOTMENTS"|"34"
360|"0454"|"CEMETERIES AND CREMATORIA"|"34"
361|"0455"|"DRINKING FOUNTAINS AND WATER POINTS"|"34"
362|"0456"|"HALLS AND COMMUNITY CENTRES"|"34"
363|"0457"|"LETTER BOXES"|"34"
364|"0458"|"LIBRARIES"|"34"
365|"0459"|"PLACES OF WORSHIP"|"34"
366|"0460"|"PUBLIC TELEPHONES"|"34"
367|"0461"|"PUBLIC TOILETS"|"34"
368|"0462"|"RECYCLING CENTRES"|"34"
369|"0802"|"WIFI HOTSPOTS"|"34"
370|"0445"|"ANIMAL WELFARE ORGANISATIONS"|"35"
371|"0446"|"FAN CLUBS AND ASSOCIATIONS"|"35"
372|"0447"|"SPORTS CLUBS AND ASSOCIATIONS"|"35"
373|"0448"|"INSTITUTES AND PROFESSIONAL ORGANISATIONS"|"35"
374|"0449"|"POLITICAL PARTIES AND RELATED ORGANISATIONS"|"35"
375|"0450"|"RELIGIOUS ORGANISATIONS"|"35"
376|"0452"|"YOUTH ORGANISATIONS"|"35"
377|"0769"|"COMMUNITY NETWORKS AND PROJECTS"|"35"
378|"0816"|"CHARITABLE ORGANISATIONS"|"35"
379|"0817"|"CONSERVATION ORGANISATIONS"|"35"
380|"0464"|"BABY, NURSERY AND PLAYGROUND EQUIPMENT"|"37"
381|"0465"|"BEDS AND BEDDING"|"37"
382|"0466"|"BRUSHES"|"37"
383|"0467"|"CANDLES"|"37"
384|"0468"|"CANVAS GOODS"|"37"
385|"0470"|"CARPETS, FLOORING, RUGS AND SOFT FURNISHINGS"|"37"
386|"0471"|"MEDALS, TROPHIES, CEREMONIAL AND RELIGIOUS GOODS"|"37"
387|"0472"|"CHINA AND GLASSWARE"|"37"
388|"0473"|"CLOTHING, COMPONENTS AND ACCESSORIES"|"37"
389|"0474"|"COOKERS AND STOVES - NON ELECTRICAL"|"37"
390|"0475"|"COSMETICS, TOILETRIES AND PERFUMES"|"37"
391|"0476"|"CURTAINS AND BLINDS"|"37"
392|"0477"|"CUTLERY AND TABLEWARE"|"37"
393|"0478"|"DISABILITY AND MOBILITY EQUIPMENT"|"37"
394|"0479"|"REFRIGERATION AND FREEZING APPLIANCES"|"37"
395|"0480"|"FOOTWEAR"|"37"
396|"0481"|"FURNITURE"|"37"
397|"0482"|"GARDEN GOODS"|"37"
398|"0483"|"GIFTWARE"|"37"
399|"0485"|"HOBBY, SPORTS AND PASTIME PRODUCTS"|"37"
400|"0486"|"DISPOSABLE PRODUCTS"|"37"
401|"0487"|"JEWELLERY, GEMS, CLOCKS AND WATCHES"|"37"
402|"0488"|"LAMPSHADES AND LIGHTING"|"37"
403|"0489"|"LEATHER PRODUCTS"|"37"
404|"0490"|"LINGERIE AND HOSIERY"|"37"
405|"0491"|"LUGGAGE, BAGS, UMBRELLAS AND TRAVEL ACCESSORIES"|"37"
406|"0493"|"MUSICAL INSTRUMENTS"|"37"
407|"0494"|"PHOTOGRAPHIC AND OPTICAL EQUIPMENT"|"37"
408|"0495"|"SAUNAS AND SUNBEDS"|"37"
409|"0497"|"TENTS, MARQUEES AND CAMPING EQUIPMENT"|"37"
410|"0498"|"TOBACCO PRODUCTS"|"37"
411|"0782"|"FIREPLACES AND MANTELPIECES"|"37"
412|"0785"|"CONSERVATORIES"|"37"
413|"0790"|"BATHROOM FIXTURES, FITTINGS AND SANITARY EQUIPMENT"|"37"
414|"0500"|"COAL MINING"|"38"
415|"0501"|"OIL AND GAS EXTRACTION, REFINERY AND PRODUCT MANUFACTURE"|"38"
416|"0502"|"ORE MINING"|"38"
417|"0503"|"PEAT EXTRACTION"|"38"
418|"0504"|"SAND, GRAVEL AND CLAY EXTRACTION AND MERCHANTS"|"38"
419|"0506"|"STONE QUARRYING AND PREPARATION"|"38"
420|"0507"|"UNSPECIFIED QUARRIES OR MINES"|"38"
421|"0508"|"ANIMAL BREEDERS (NOT HORSES)"|"39"
422|"0509"|"ARABLE FARMING"|"39"
423|"0510"|"BEE KEEPERS"|"39"
424|"0511"|"DAIRY FARMING"|"39"
425|"0512"|"FISH AND SHELLFISH"|"39"
426|"0513"|"FORESTRY"|"39"
427|"0514"|"FRUIT, FLOWER AND VEGETABLE GROWERS"|"39"
428|"0515"|"HOPPERS AND SILOS"|"39"
429|"0516"|"HORSE BREEDERS AND DEALERS"|"39"
430|"0517"|"LIVESTOCK FARMING"|"39"
431|"0518"|"MIXED OR UNSPECIFIED FARMING"|"39"
432|"0520"|"POULTRY FARMING, EQUIPMENT AND SUPPLIES"|"39"
433|"0521"|"SHEEP DIPS AND WASHES"|"39"
434|"0522"|"ALCOHOLIC DRINKS"|"40"
435|"0523"|"ANIMAL FEEDS, PET FOODS, HAY AND STRAW"|"40"
436|"0524"|"BAKING AND CONFECTIONERY"|"40"
437|"0525"|"DAIRY PRODUCTS"|"40"
438|"0526"|"FISH, MEAT AND POULTRY PRODUCTS"|"40"
439|"0528"|"MILLING, REFINING AND FOOD ADDITIVES"|"40"
440|"0529"|"NON ALCOHOLIC DRINKS"|"40"
441|"0530"|"CATERING AND NON SPECIFIC FOOD PRODUCTS"|"40"
442|"0531"|"BUSINESS PARKS AND INDUSTRIAL ESTATES"|"41"
443|"0532"|"CHIMNEYS"|"41"
444|"0533"|"CONVEYORS"|"41"
445|"0534"|"ENERGY PRODUCTION"|"41"
446|"0535"|"LIGHTING TOWERS"|"41"
447|"0536"|"LIME KILNS"|"41"
448|"0537"|"OAST HOUSES"|"41"
449|"0538"|"PIPELINES"|"41"
450|"0539"|"TANKS (GENERIC)"|"41"
451|"0540"|"TRAVELLING CRANES AND GANTRIES"|"41"
452|"0542"|"UNSPECIFIED WORKS OR FACTORIES"|"41"
453|"0543"|"WATER PUMPING STATIONS"|"41"
454|"0544"|"ABRASIVE PRODUCTS AND GRINDING EQUIPMENT"|"42"
455|"0545"|"ADHESIVES AND SEALANTS"|"42"
456|"0546"|"AEROPLANES"|"42"
457|"0547"|"AGRICULTURAL MACHINERY AND GOODS"|"42"
458|"0548"|"AIR AND WATER FILTRATION"|"42"
459|"0549"|"ARMS AND AMMUNITION"|"42"
460|"0550"|"BEARING, GEAR AND DRIVE ELEMENTS"|"42"
461|"0551"|"BEEKEEPING SUPPLIES"|"42"
462|"0553"|"BRICKS, TILES, CLAY AND CERAMIC PRODUCTS"|"42"
463|"0555"|"CABLE, WIRE AND FIBRE OPTICS"|"42"
464|"0557"|"COLOURS, CHEMICALS AND WATER SOFTENERS AND SUPPLIES"|"42"
465|"0558"|"CLEANING EQUIPMENT AND SUPPLIES"|"42"
466|"0562"|"CONCRETE PRODUCTS"|"42"
467|"0563"|"COOLING AND REFRIGERATION"|"42"
468|"0564"|"ELECTRICAL COMPONENTS"|"42"
469|"0565"|"ELECTRICAL MOTORS AND GENERATORS"|"42"
470|"0566"|"ELECTRICAL PRODUCTION AND MANIPULATION EQUIPMENT"|"42"
471|"0567"|"ELECTRONIC EQUIPMENT"|"42"
472|"0568"|"ELECTRONIC MEDIA"|"42"
473|"0569"|"ENGINES"|"42"
474|"0571"|"FERTILISERS"|"42"
475|"0572"|"FOOD AND BEVERAGE INDUSTRY MACHINERY"|"42"
476|"0573"|"GENERAL CONSTRUCTION SUPPLIES"|"42"
477|"0574"|"GENERAL PURPOSE MACHINERY"|"42"
478|"0575"|"GLASS"|"42"
479|"0576"|"HORTICULTURAL EQUIPMENT"|"42"
480|"0577"|"INDUSTRIAL COATINGS AND FINISHINGS"|"42"
481|"0579"|"TOOLS INCLUDING MACHINE SHOPS"|"42"
482|"0580"|"LIFTING AND HANDLING EQUIPMENT"|"42"
483|"0581"|"LUBRICANTS AND LUBRICATING EQUIPMENT"|"42"
484|"0582"|"MARINE EQUIPMENT INCLUDING BOATS AND SHIPS"|"42"
485|"0583"|"MEASUREMENT AND INSPECTION EQUIPMENT"|"42"
486|"0584"|"MEDICAL EQUIPMENT, SUPPLIES AND PHARMACEUTICALS"|"42"
487|"0585"|"METALS MANUFACTURERS, FABRICATORS AND STOCKHOLDERS"|"42"
488|"0586"|"MOULDS, DIES AND CASTINGS"|"42"
489|"0588"|"OFFICE AND SHOP EQUIPMENT"|"42"
490|"0589"|"OVENS AND FURNACES"|"42"
491|"0590"|"PACKAGING"|"42"
492|"0591"|"PAINTS, VARNISHES AND LACQUERS"|"42"
493|"0594"|"PESTICIDES"|"42"
494|"0598"|"PRINTING RELATED MACHINERY"|"42"
495|"0599"|"PUBLISHED GOODS"|"42"
496|"0600"|"PUMPS AND COMPRESSORS"|"42"
497|"0601"|"RADAR AND TELECOMMUNICATIONS EQUIPMENT"|"42"
498|"0602"|"ROAD MAINTENANCE EQUIPMENT"|"42"
499|"0603"|"ROPES, NETS AND CORDAGE"|"42"
500|"0604"|"RUBBER, SILICONES AND PLASTICS"|"42"
501|"0605"|"SEALS, TAPES, TAPS AND VALVES"|"42"
502|"0606"|"SIGNS"|"42"
503|"0607"|"SPECIAL PURPOSE MACHINERY AND EQUIPMENT"|"42"
504|"0608"|"TEXTILES, FABRICS, SILK AND MACHINERY"|"42"
505|"0609"|"STATIONERY, STAMPS, TAGS AND LABELS"|"42"
506|"0612"|"GENERAL MANUFACTURING"|"42"
507|"0613"|"VEHICLE BODYBUILDERS"|"42"
508|"0614"|"VEHICLE COMPONENTS"|"42"
509|"0615"|"VEHICLES"|"42"
510|"0616"|"WOOD PRODUCTS INCLUDING CHARCOAL, PAPER, CARD AND BOARD"|"42"
511|"0617"|"WORKWEAR"|"42"
512|"0765"|"EDUCATIONAL EQUIPMENT AND SUPPLIES"|"42"
513|"0767"|"ICE"|"42"
514|"0781"|"FENCES, GATES AND RAILINGS"|"42"
515|"0783"|"ACCESS EQUIPMENT"|"42"
516|"0784"|"CAR PORTS AND STEEL BUILDINGS"|"42"
517|"0787"|"WASTE COLLECTION, PROCESSING AND DISPOSAL EQUIPMENT"|"42"
518|"0788"|"GLASS FIBRE SERVICES"|"42"
519|"0791"|"SHELVING, STORAGE, SAFES AND VAULTS"|"42"
520|"0656"|"CLOTHING"|"46"
521|"0657"|"FOOTWEAR"|"46"
522|"0659"|"JEWELLERY AND FASHION ACCESSORIES"|"46"
523|"0660"|"LINGERIE AND HOSIERY"|"46"
524|"0797"|"BABY AND NURSERY EQUIPMENT AND CHILDREN'S CLOTHES"|"46"
525|"0661"|"BAKERIES"|"47"
526|"0662"|"BUTCHERS"|"47"
527|"0663"|"CONFECTIONERS"|"47"
528|"0665"|"DELICATESSENS"|"47"
529|"0666"|"FISHMONGERS"|"47"
530|"0667"|"FROZEN FOODS"|"47"
531|"0668"|"GREEN AND NEW AGE GOODS"|"47"
532|"0669"|"GROCERS, FARM SHOPS AND PICK YOUR OWN"|"47"
533|"0670"|"HERBS AND SPICES"|"47"
534|"0671"|"ALCOHOLIC DRINKS INCLUDING OFF LICENCES AND WHOLESALERS"|"47"
535|"0672"|"ORGANIC, HEALTH, GOURMET AND KOSHER FOODS"|"47"
536|"0699"|"CONVENIENCE STORES AND INDEPENDENT SUPERMARKETS"|"47"
537|"0703"|"LIVESTOCK MARKETS"|"47"
538|"0705"|"MARKETS"|"47"
539|"0768"|"CASH AND CARRY"|"47"
540|"0798"|"TEA AND COFFEE MERCHANTS"|"47"
541|"0819"|"SUPERMARKET CHAINS"|"47"
542|"0674"|"BOOKS AND MAPS"|"48"
543|"0675"|"CARPETS, RUGS, SOFT FURNISHINGS AND NEEDLECRAFT"|"48"
544|"0676"|"CHINA AND GLASSWARE"|"48"
545|"0677"|"COSMETICS, TOILETRIES, PERFUMES AND HAIRDRESSING SUPPLIES"|"48"
546|"0678"|"CRAFT SUPPLIES"|"48"
547|"0679"|"CYCLES AND ACCESSORIES"|"48"
548|"0680"|"DIY AND HOME IMPROVEMENT"|"48"
549|"0682"|"FURNITURE"|"48"
550|"0683"|"GARDEN CENTRES AND NURSERIES"|"48"
551|"0684"|"GARDEN MACHINERY AND FURNITURE"|"48"
552|"0685"|"GENERAL HOUSEHOLD GOODS"|"48"
553|"0686"|"HOBBY, SPORTS AND PASTIME PRODUCTS"|"48"
554|"0687"|"LEATHER GOODS, LUGGAGE AND TRAVEL ACCESSORIES INCLUDING HANDBAGS"|"48"
555|"0688"|"LIGHTING"|"48"
556|"0689"|"MUSIC AND VIDEO"|"48"
557|"0690"|"MUSICAL INSTRUMENTS"|"48"
558|"0691"|"PETS, SUPPLIES AND SERVICES"|"48"
559|"0693"|"CAMPING AND CARAVANNING"|"48"
560|"0694"|"TRAVEL AGENCIES"|"48"
561|"0700"|"DEPARTMENT STORES"|"48"
562|"0701"|"DISCOUNT STORES"|"48"
563|"0704"|"MAIL ORDER AND CATALOGUE STORES"|"48"
564|"0708"|"SHOPPING CENTRES AND RETAIL PARKS"|"48"
565|"0710"|"SURPLUS GOODS"|"48"
566|"0712"|"ART AND ANTIQUES"|"48"
567|"0714"|"CHARITY SHOPS"|"48"
568|"0716"|"FLORISTS"|"48"
569|"0717"|"GIFTS AND CARDS"|"48"
570|"0718"|"PARTY GOODS AND NOVELTIES"|"48"
571|"0719"|"SECONDHAND GOODS"|"48"
572|"0720"|"COMPUTER SUPPLIES"|"48"
573|"0721"|"DOMESTIC APPLIANCES"|"48"
574|"0722"|"ELECTRICAL GOODS AND COMPONENTS"|"48"
575|"0724"|"PHOTOGRAPHIC AND OPTICAL EQUIPMENT"|"48"
576|"0725"|"STATIONERY AND OFFICE SUPPLIES"|"48"
577|"0726"|"TELEPHONES AND TELEPHONE CARDS"|"48"
578|"0763"|"POST OFFICES"|"48"
579|"0764"|"GARAGES, GARDEN AND PORTABLE BUILDINGS"|"48"
580|"0766"|"FUEL DISTRIBUTORS AND SUPPLIERS"|"48"
581|"0824"|"ADULT SHOPS"|"48"
582|"0827"|"COMICS BOOKSHOPS"|"48"
583|"0828"|"COMPUTER SHOPS"|"48"
584|"0831"|"POTTERIES"|"48"
585|"0695"|"NEW VEHICLES"|"49"
586|"0696"|"SECONDHAND VEHICLES"|"49"
587|"0697"|"VEHICLE AUCTIONS"|"49"
588|"0698"|"VEHICLE PARTS AND ACCESSORIES"|"49"
589|"0727"|"AERONAUTICAL FEATURES"|"53"
590|"0728"|"AIRPORTS AND LANDING STRIPS"|"53"
591|"0729"|"HELIPADS"|"53"
592|"0730"|"BRIDGES"|"54"
593|"0733"|"CATTLE GRIDS"|"54"
594|"0734"|"FORDS AND LEVEL CROSSINGS"|"54"
595|"0735"|"MOTORWAY SERVICE STATIONS"|"54"
596|"0736"|"PARKING"|"54"
597|"0737"|"PETROL AND FUEL STATIONS"|"54"
598|"0739"|"ROADSIDE TELEPHONE BOXES"|"54"
599|"0740"|"SIGNALLING FACILITIES"|"54"
600|"0742"|"TUNNELS"|"54"
601|"0743"|"VIADUCTS"|"54"
602|"0744"|"WEIGHBRIDGES"|"54"
603|"0746"|"FINGER POSTS, GUIDE POSTS AND CAIRNS"|"55"
604|"0747"|"FOOTBRIDGES"|"55"
605|"0749"|"STEPPING STONES"|"55"
606|"0750"|"SUBWAYS"|"55"
607|"0751"|"AQUEDUCTS"|"56"
608|"0752"|"LOCKS"|"56"
609|"0753"|"MOORINGS AND UNLOADING FACILITIES"|"56"
610|"0754"|"RIVERS AND CANAL ORGANISATIONS AND INFRASTRUCTURE"|"56"
611|"0755"|"WEIRS, SLUICES AND DAMS"|"56"
612|"0760"|"FERRIES AND FERRY TERMINALS"|"56"
613|"0731"|"BUS AND COACH STATIONS, DEPOTS AND COMPANIES"|"57"
614|"0738"|"RAILWAY STATIONS, JUNCTIONS AND HALTS"|"57"
615|"0756"|"TRAM, METRO AND LIGHT RAILWAY STATIONS AND STOPS"|"57"
616|"0758"|"TAXI RANKS"|"57"
617|"0761"|"UNDERGROUND NETWORK STATIONS"|"57"
618|"0794"|"LONDON UNDERGROUND ENTRANCES"|"57"
619|"0732"|"BUS STOPS"|"59"
620|"0759"|"HAIL AND RIDE ZONES"|"59"
